module Calculator(
    input [31:0] addra,
    input [7:0] ascii_in,
    input [15:0] kbsig,//8:u, 7:d, 6:l, 5:r
    input clk,
    input in_valid,
    output [11:0] douta,
    input available
);
    wire out;
    reg [7:0] text [2399:0];
    reg [31:0] ptr = 80;
    initial begin
        text[0] = 8'd84;
        text[1] = 8'd66;
        text[2] = 8'd68;
        text[3] = 8'd0;
        text[4] = 8'd0;
        text[5] = 8'd0;
        text[6] = 8'd0;
        text[7] = 8'd0;
        text[8] = 8'd0;
        text[9] = 8'd0;
        text[10] = 8'd0;
        text[11] = 8'd0;
        text[12] = 8'd0;
        text[13] = 8'd0;
        text[14] = 8'd0;
        text[15] = 8'd0;
        text[16] = 8'd0;
        text[17] = 8'd0;
        text[18] = 8'd0;
        text[19] = 8'd0;
        text[20] = 8'd0;
        text[21] = 8'd0;
        text[22] = 8'd0;
        text[23] = 8'd0;
        text[24] = 8'd0;
        text[25] = 8'd0;
        text[26] = 8'd0;
        text[27] = 8'd0;
        text[28] = 8'd0;
        text[29] = 8'd0;
        text[30] = 8'd0;
        text[31] = 8'd0;
        text[32] = 8'd0;
        text[33] = 8'd0;
        text[34] = 8'd0;
        text[35] = 8'd0;
        text[36] = 8'd0;
        text[37] = 8'd0;
        text[38] = 8'd0;
        text[39] = 8'd0;
        text[40] = 8'd0;
        text[41] = 8'd0;
        text[42] = 8'd0;
        text[43] = 8'd0;
        text[44] = 8'd0;
        text[45] = 8'd0;
        text[46] = 8'd0;
        text[47] = 8'd0;
        text[48] = 8'd0;
        text[49] = 8'd0;
        text[50] = 8'd0;
        text[51] = 8'd0;
        text[52] = 8'd0;
        text[53] = 8'd0;
        text[54] = 8'd0;
        text[55] = 8'd0;
        text[56] = 8'd0;
        text[57] = 8'd0;
        text[58] = 8'd0;
        text[59] = 8'd0;
        text[60] = 8'd0;
        text[61] = 8'd0;
        text[62] = 8'd0;
        text[63] = 8'd0;
        text[64] = 8'd0;
        text[65] = 8'd0;
        text[66] = 8'd0;
        text[67] = 8'd0;
        text[68] = 8'd0;
        text[69] = 8'd0;
        text[70] = 8'd0;
        text[71] = 8'd0;
        text[72] = 8'd0;
        text[73] = 8'd0;
        text[74] = 8'd0;
        text[75] = 8'd0;
        text[76] = 8'd0;
        text[77] = 8'd0;
        text[78] = 8'd0;
        text[79] = 8'd0;
        text[80] = 8'd73;
        text[81] = 8'd39;
        text[82] = 8'd118;
        text[83] = 8'd101;
        text[84] = 8'd32;
        text[85] = 8'd103;
        text[86] = 8'd111;
        text[87] = 8'd116;
        text[88] = 8'd32;
        text[89] = 8'd115;
        text[90] = 8'd111;
        text[91] = 8'd109;
        text[92] = 8'd101;
        text[93] = 8'd32;
        text[94] = 8'd104;
        text[95] = 8'd111;
        text[96] = 8'd116;
        text[97] = 8'd32;
        text[98] = 8'd112;
        text[99] = 8'd111;
        text[100] = 8'd116;
        text[101] = 8'd97;
        text[102] = 8'd116;
        text[103] = 8'd111;
        text[104] = 8'd101;
        text[105] = 8'd115;
        text[106] = 8'd32;
        text[107] = 8'd111;
        text[108] = 8'd110;
        text[109] = 8'd32;
        text[110] = 8'd109;
        text[111] = 8'd121;
        text[112] = 8'd32;
        text[113] = 8'd104;
        text[114] = 8'd97;
        text[115] = 8'd110;
        text[116] = 8'd100;
        text[117] = 8'd115;
        text[118] = 8'd46;
        text[119] = 8'd0;
        text[120] = 8'd0;
        text[121] = 8'd0;
        text[122] = 8'd0;
        text[123] = 8'd0;
        text[124] = 8'd0;
        text[125] = 8'd0;
        text[126] = 8'd0;
        text[127] = 8'd0;
        text[128] = 8'd0;
        text[129] = 8'd0;
        text[130] = 8'd0;
        text[131] = 8'd0;
        text[132] = 8'd0;
        text[133] = 8'd0;
        text[134] = 8'd0;
        text[135] = 8'd0;
        text[136] = 8'd0;
        text[137] = 8'd0;
        text[138] = 8'd0;
        text[139] = 8'd0;
        text[140] = 8'd0;
        text[141] = 8'd0;
        text[142] = 8'd0;
        text[143] = 8'd0;
        text[144] = 8'd0;
        text[145] = 8'd0;
        text[146] = 8'd0;
        text[147] = 8'd0;
        text[148] = 8'd0;
        text[149] = 8'd0;
        text[150] = 8'd0;
        text[151] = 8'd0;
        text[152] = 8'd0;
        text[153] = 8'd0;
        text[154] = 8'd0;
        text[155] = 8'd0;
        text[156] = 8'd0;
        text[157] = 8'd0;
        text[158] = 8'd0;
        text[159] = 8'd0;
    end
    wire [31:0] xw = addra % 8, yw = ((addra / 640) % 16);
    wire [31:0] caddr;
    assign caddr = 80 * (addra / (640 * 16)) + (((addra % (640 * 16)) / 8) % 80);
    get_charpix pix(
        .c(caddr >= 160 ? 0 : text[caddr]),
        .x(xw[5:0]),
        .y(yw[5:0]),
        .in_ptr((80 * (addra / (640 * 16)) + (((addra % (640 * 16)) / 8) % 80)) == ptr),
        .is_light(out)
    );
    assign douta = (out == 1) ? 12'b111111111111 : 12'd0; 
endmodule