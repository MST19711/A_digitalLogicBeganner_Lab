`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/10/02 00:39:53
// Design Name: 
// Module Name: mul_32p
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module adder_1(
    input a,
    input b,
    input cin,
    output f,
    output cout
);
    assign f = (a ^ b) ^ cin;
    assign cout =  (a & b) | (a & cin) | (b & cin);
endmodule

module mul_32k(
    input [31:0] X, Y,
    output reg [63:0] P       // output variable for assignment
);
//add your code here  
    wire [31:0] L0;
    wire [31:0] C0 = 32'b0;
    /*
    ```python3
        for i in range(0, 32):
            print("assign L0[{}] = X[{}] & Y[0];".format(str(i), str(i)))
    ```
    */
    assign L0[0] = X[0] & Y[0];
    assign L0[1] = X[1] & Y[0];
    assign L0[2] = X[2] & Y[0];
    assign L0[3] = X[3] & Y[0];
    assign L0[4] = X[4] & Y[0];
    assign L0[5] = X[5] & Y[0];
    assign L0[6] = X[6] & Y[0];
    assign L0[7] = X[7] & Y[0];
    assign L0[8] = X[8] & Y[0];
    assign L0[9] = X[9] & Y[0];
    assign L0[10] = X[10] & Y[0];
    assign L0[11] = X[11] & Y[0];
    assign L0[12] = X[12] & Y[0];
    assign L0[13] = X[13] & Y[0];
    assign L0[14] = X[14] & Y[0];
    assign L0[15] = X[15] & Y[0];
    assign L0[16] = X[16] & Y[0];
    assign L0[17] = X[17] & Y[0];
    assign L0[18] = X[18] & Y[0];
    assign L0[19] = X[19] & Y[0];
    assign L0[20] = X[20] & Y[0];
    assign L0[21] = X[21] & Y[0];
    assign L0[22] = X[22] & Y[0];
    assign L0[23] = X[23] & Y[0];
    assign L0[24] = X[24] & Y[0];
    assign L0[25] = X[25] & Y[0];
    assign L0[26] = X[26] & Y[0];
    assign L0[27] = X[27] & Y[0];
    assign L0[28] = X[28] & Y[0];
    assign L0[29] = X[29] & Y[0];
    assign L0[30] = X[30] & Y[0];
    assign L0[31] = X[31] & Y[0];
    /*
    ```python3
        for i in range(1, 32):
            print("wire [31:0] L{}, C{};".format(str(i), str(i)))
            for j in range(0, 31):
                print("adder_1 adder{}(.a(X[{}] & Y[{}]), .b(L{}[{}]), .cin(C{}[{}]), .f(L{}[{}]), .cout(C{}[{}]));".format(str(i) + "_" + str(j), str(j), str(i), str(i-1), str(j+1), str(i-1), str(j), str(i), str(j), str(i), str(j)))
            print("assign L{}[31] = X[31] & Y[{}];".format(str(i), str(i)))
            print("assign P[{}] = L{}[0];".format(str(i), str(i)))
    ```
    */
    wire [31:0] L1, C1;
    adder_1 adder1_0(.a(X[0] & Y[1]), .b(L0[1]), .cin(C0[0]), .f(L1[0]), .cout(C1[0]));
    adder_1 adder1_1(.a(X[1] & Y[1]), .b(L0[2]), .cin(C0[1]), .f(L1[1]), .cout(C1[1]));
    adder_1 adder1_2(.a(X[2] & Y[1]), .b(L0[3]), .cin(C0[2]), .f(L1[2]), .cout(C1[2]));
    adder_1 adder1_3(.a(X[3] & Y[1]), .b(L0[4]), .cin(C0[3]), .f(L1[3]), .cout(C1[3]));
    adder_1 adder1_4(.a(X[4] & Y[1]), .b(L0[5]), .cin(C0[4]), .f(L1[4]), .cout(C1[4]));
    adder_1 adder1_5(.a(X[5] & Y[1]), .b(L0[6]), .cin(C0[5]), .f(L1[5]), .cout(C1[5]));
    adder_1 adder1_6(.a(X[6] & Y[1]), .b(L0[7]), .cin(C0[6]), .f(L1[6]), .cout(C1[6]));
    adder_1 adder1_7(.a(X[7] & Y[1]), .b(L0[8]), .cin(C0[7]), .f(L1[7]), .cout(C1[7]));
    adder_1 adder1_8(.a(X[8] & Y[1]), .b(L0[9]), .cin(C0[8]), .f(L1[8]), .cout(C1[8]));
    adder_1 adder1_9(.a(X[9] & Y[1]), .b(L0[10]), .cin(C0[9]), .f(L1[9]), .cout(C1[9]));
    adder_1 adder1_10(.a(X[10] & Y[1]), .b(L0[11]), .cin(C0[10]), .f(L1[10]), .cout(C1[10]));
    adder_1 adder1_11(.a(X[11] & Y[1]), .b(L0[12]), .cin(C0[11]), .f(L1[11]), .cout(C1[11]));
    adder_1 adder1_12(.a(X[12] & Y[1]), .b(L0[13]), .cin(C0[12]), .f(L1[12]), .cout(C1[12]));
    adder_1 adder1_13(.a(X[13] & Y[1]), .b(L0[14]), .cin(C0[13]), .f(L1[13]), .cout(C1[13]));
    adder_1 adder1_14(.a(X[14] & Y[1]), .b(L0[15]), .cin(C0[14]), .f(L1[14]), .cout(C1[14]));
    adder_1 adder1_15(.a(X[15] & Y[1]), .b(L0[16]), .cin(C0[15]), .f(L1[15]), .cout(C1[15]));
    adder_1 adder1_16(.a(X[16] & Y[1]), .b(L0[17]), .cin(C0[16]), .f(L1[16]), .cout(C1[16]));
    adder_1 adder1_17(.a(X[17] & Y[1]), .b(L0[18]), .cin(C0[17]), .f(L1[17]), .cout(C1[17]));
    adder_1 adder1_18(.a(X[18] & Y[1]), .b(L0[19]), .cin(C0[18]), .f(L1[18]), .cout(C1[18]));
    adder_1 adder1_19(.a(X[19] & Y[1]), .b(L0[20]), .cin(C0[19]), .f(L1[19]), .cout(C1[19]));
    adder_1 adder1_20(.a(X[20] & Y[1]), .b(L0[21]), .cin(C0[20]), .f(L1[20]), .cout(C1[20]));
    adder_1 adder1_21(.a(X[21] & Y[1]), .b(L0[22]), .cin(C0[21]), .f(L1[21]), .cout(C1[21]));
    adder_1 adder1_22(.a(X[22] & Y[1]), .b(L0[23]), .cin(C0[22]), .f(L1[22]), .cout(C1[22]));
    adder_1 adder1_23(.a(X[23] & Y[1]), .b(L0[24]), .cin(C0[23]), .f(L1[23]), .cout(C1[23]));
    adder_1 adder1_24(.a(X[24] & Y[1]), .b(L0[25]), .cin(C0[24]), .f(L1[24]), .cout(C1[24]));
    adder_1 adder1_25(.a(X[25] & Y[1]), .b(L0[26]), .cin(C0[25]), .f(L1[25]), .cout(C1[25]));
    adder_1 adder1_26(.a(X[26] & Y[1]), .b(L0[27]), .cin(C0[26]), .f(L1[26]), .cout(C1[26]));
    adder_1 adder1_27(.a(X[27] & Y[1]), .b(L0[28]), .cin(C0[27]), .f(L1[27]), .cout(C1[27]));
    adder_1 adder1_28(.a(X[28] & Y[1]), .b(L0[29]), .cin(C0[28]), .f(L1[28]), .cout(C1[28]));
    adder_1 adder1_29(.a(X[29] & Y[1]), .b(L0[30]), .cin(C0[29]), .f(L1[29]), .cout(C1[29]));
    adder_1 adder1_30(.a(X[30] & Y[1]), .b(L0[31]), .cin(C0[30]), .f(L1[30]), .cout(C1[30]));
    assign L1[31] = X[31] & Y[1];
    wire [31:0] L2, C2;
    adder_1 adder2_0(.a(X[0] & Y[2]), .b(L1[1]), .cin(C1[0]), .f(L2[0]), .cout(C2[0]));
    adder_1 adder2_1(.a(X[1] & Y[2]), .b(L1[2]), .cin(C1[1]), .f(L2[1]), .cout(C2[1]));
    adder_1 adder2_2(.a(X[2] & Y[2]), .b(L1[3]), .cin(C1[2]), .f(L2[2]), .cout(C2[2]));
    adder_1 adder2_3(.a(X[3] & Y[2]), .b(L1[4]), .cin(C1[3]), .f(L2[3]), .cout(C2[3]));
    adder_1 adder2_4(.a(X[4] & Y[2]), .b(L1[5]), .cin(C1[4]), .f(L2[4]), .cout(C2[4]));
    adder_1 adder2_5(.a(X[5] & Y[2]), .b(L1[6]), .cin(C1[5]), .f(L2[5]), .cout(C2[5]));
    adder_1 adder2_6(.a(X[6] & Y[2]), .b(L1[7]), .cin(C1[6]), .f(L2[6]), .cout(C2[6]));
    adder_1 adder2_7(.a(X[7] & Y[2]), .b(L1[8]), .cin(C1[7]), .f(L2[7]), .cout(C2[7]));
    adder_1 adder2_8(.a(X[8] & Y[2]), .b(L1[9]), .cin(C1[8]), .f(L2[8]), .cout(C2[8]));
    adder_1 adder2_9(.a(X[9] & Y[2]), .b(L1[10]), .cin(C1[9]), .f(L2[9]), .cout(C2[9]));
    adder_1 adder2_10(.a(X[10] & Y[2]), .b(L1[11]), .cin(C1[10]), .f(L2[10]), .cout(C2[10]));
    adder_1 adder2_11(.a(X[11] & Y[2]), .b(L1[12]), .cin(C1[11]), .f(L2[11]), .cout(C2[11]));
    adder_1 adder2_12(.a(X[12] & Y[2]), .b(L1[13]), .cin(C1[12]), .f(L2[12]), .cout(C2[12]));
    adder_1 adder2_13(.a(X[13] & Y[2]), .b(L1[14]), .cin(C1[13]), .f(L2[13]), .cout(C2[13]));
    adder_1 adder2_14(.a(X[14] & Y[2]), .b(L1[15]), .cin(C1[14]), .f(L2[14]), .cout(C2[14]));
    adder_1 adder2_15(.a(X[15] & Y[2]), .b(L1[16]), .cin(C1[15]), .f(L2[15]), .cout(C2[15]));
    adder_1 adder2_16(.a(X[16] & Y[2]), .b(L1[17]), .cin(C1[16]), .f(L2[16]), .cout(C2[16]));
    adder_1 adder2_17(.a(X[17] & Y[2]), .b(L1[18]), .cin(C1[17]), .f(L2[17]), .cout(C2[17]));
    adder_1 adder2_18(.a(X[18] & Y[2]), .b(L1[19]), .cin(C1[18]), .f(L2[18]), .cout(C2[18]));
    adder_1 adder2_19(.a(X[19] & Y[2]), .b(L1[20]), .cin(C1[19]), .f(L2[19]), .cout(C2[19]));
    adder_1 adder2_20(.a(X[20] & Y[2]), .b(L1[21]), .cin(C1[20]), .f(L2[20]), .cout(C2[20]));
    adder_1 adder2_21(.a(X[21] & Y[2]), .b(L1[22]), .cin(C1[21]), .f(L2[21]), .cout(C2[21]));
    adder_1 adder2_22(.a(X[22] & Y[2]), .b(L1[23]), .cin(C1[22]), .f(L2[22]), .cout(C2[22]));
    adder_1 adder2_23(.a(X[23] & Y[2]), .b(L1[24]), .cin(C1[23]), .f(L2[23]), .cout(C2[23]));
    adder_1 adder2_24(.a(X[24] & Y[2]), .b(L1[25]), .cin(C1[24]), .f(L2[24]), .cout(C2[24]));
    adder_1 adder2_25(.a(X[25] & Y[2]), .b(L1[26]), .cin(C1[25]), .f(L2[25]), .cout(C2[25]));
    adder_1 adder2_26(.a(X[26] & Y[2]), .b(L1[27]), .cin(C1[26]), .f(L2[26]), .cout(C2[26]));
    adder_1 adder2_27(.a(X[27] & Y[2]), .b(L1[28]), .cin(C1[27]), .f(L2[27]), .cout(C2[27]));
    adder_1 adder2_28(.a(X[28] & Y[2]), .b(L1[29]), .cin(C1[28]), .f(L2[28]), .cout(C2[28]));
    adder_1 adder2_29(.a(X[29] & Y[2]), .b(L1[30]), .cin(C1[29]), .f(L2[29]), .cout(C2[29]));
    adder_1 adder2_30(.a(X[30] & Y[2]), .b(L1[31]), .cin(C1[30]), .f(L2[30]), .cout(C2[30]));
    assign L2[31] = X[31] & Y[2];
    wire [31:0] L3, C3;
    adder_1 adder3_0(.a(X[0] & Y[3]), .b(L2[1]), .cin(C2[0]), .f(L3[0]), .cout(C3[0]));
    adder_1 adder3_1(.a(X[1] & Y[3]), .b(L2[2]), .cin(C2[1]), .f(L3[1]), .cout(C3[1]));
    adder_1 adder3_2(.a(X[2] & Y[3]), .b(L2[3]), .cin(C2[2]), .f(L3[2]), .cout(C3[2]));
    adder_1 adder3_3(.a(X[3] & Y[3]), .b(L2[4]), .cin(C2[3]), .f(L3[3]), .cout(C3[3]));
    adder_1 adder3_4(.a(X[4] & Y[3]), .b(L2[5]), .cin(C2[4]), .f(L3[4]), .cout(C3[4]));
    adder_1 adder3_5(.a(X[5] & Y[3]), .b(L2[6]), .cin(C2[5]), .f(L3[5]), .cout(C3[5]));
    adder_1 adder3_6(.a(X[6] & Y[3]), .b(L2[7]), .cin(C2[6]), .f(L3[6]), .cout(C3[6]));
    adder_1 adder3_7(.a(X[7] & Y[3]), .b(L2[8]), .cin(C2[7]), .f(L3[7]), .cout(C3[7]));
    adder_1 adder3_8(.a(X[8] & Y[3]), .b(L2[9]), .cin(C2[8]), .f(L3[8]), .cout(C3[8]));
    adder_1 adder3_9(.a(X[9] & Y[3]), .b(L2[10]), .cin(C2[9]), .f(L3[9]), .cout(C3[9]));
    adder_1 adder3_10(.a(X[10] & Y[3]), .b(L2[11]), .cin(C2[10]), .f(L3[10]), .cout(C3[10]));
    adder_1 adder3_11(.a(X[11] & Y[3]), .b(L2[12]), .cin(C2[11]), .f(L3[11]), .cout(C3[11]));
    adder_1 adder3_12(.a(X[12] & Y[3]), .b(L2[13]), .cin(C2[12]), .f(L3[12]), .cout(C3[12]));
    adder_1 adder3_13(.a(X[13] & Y[3]), .b(L2[14]), .cin(C2[13]), .f(L3[13]), .cout(C3[13]));
    adder_1 adder3_14(.a(X[14] & Y[3]), .b(L2[15]), .cin(C2[14]), .f(L3[14]), .cout(C3[14]));
    adder_1 adder3_15(.a(X[15] & Y[3]), .b(L2[16]), .cin(C2[15]), .f(L3[15]), .cout(C3[15]));
    adder_1 adder3_16(.a(X[16] & Y[3]), .b(L2[17]), .cin(C2[16]), .f(L3[16]), .cout(C3[16]));
    adder_1 adder3_17(.a(X[17] & Y[3]), .b(L2[18]), .cin(C2[17]), .f(L3[17]), .cout(C3[17]));
    adder_1 adder3_18(.a(X[18] & Y[3]), .b(L2[19]), .cin(C2[18]), .f(L3[18]), .cout(C3[18]));
    adder_1 adder3_19(.a(X[19] & Y[3]), .b(L2[20]), .cin(C2[19]), .f(L3[19]), .cout(C3[19]));
    adder_1 adder3_20(.a(X[20] & Y[3]), .b(L2[21]), .cin(C2[20]), .f(L3[20]), .cout(C3[20]));
    adder_1 adder3_21(.a(X[21] & Y[3]), .b(L2[22]), .cin(C2[21]), .f(L3[21]), .cout(C3[21]));
    adder_1 adder3_22(.a(X[22] & Y[3]), .b(L2[23]), .cin(C2[22]), .f(L3[22]), .cout(C3[22]));
    adder_1 adder3_23(.a(X[23] & Y[3]), .b(L2[24]), .cin(C2[23]), .f(L3[23]), .cout(C3[23]));
    adder_1 adder3_24(.a(X[24] & Y[3]), .b(L2[25]), .cin(C2[24]), .f(L3[24]), .cout(C3[24]));
    adder_1 adder3_25(.a(X[25] & Y[3]), .b(L2[26]), .cin(C2[25]), .f(L3[25]), .cout(C3[25]));
    adder_1 adder3_26(.a(X[26] & Y[3]), .b(L2[27]), .cin(C2[26]), .f(L3[26]), .cout(C3[26]));
    adder_1 adder3_27(.a(X[27] & Y[3]), .b(L2[28]), .cin(C2[27]), .f(L3[27]), .cout(C3[27]));
    adder_1 adder3_28(.a(X[28] & Y[3]), .b(L2[29]), .cin(C2[28]), .f(L3[28]), .cout(C3[28]));
    adder_1 adder3_29(.a(X[29] & Y[3]), .b(L2[30]), .cin(C2[29]), .f(L3[29]), .cout(C3[29]));
    adder_1 adder3_30(.a(X[30] & Y[3]), .b(L2[31]), .cin(C2[30]), .f(L3[30]), .cout(C3[30]));
    assign L3[31] = X[31] & Y[3];
    wire [31:0] L4, C4;
    adder_1 adder4_0(.a(X[0] & Y[4]), .b(L3[1]), .cin(C3[0]), .f(L4[0]), .cout(C4[0]));
    adder_1 adder4_1(.a(X[1] & Y[4]), .b(L3[2]), .cin(C3[1]), .f(L4[1]), .cout(C4[1]));
    adder_1 adder4_2(.a(X[2] & Y[4]), .b(L3[3]), .cin(C3[2]), .f(L4[2]), .cout(C4[2]));
    adder_1 adder4_3(.a(X[3] & Y[4]), .b(L3[4]), .cin(C3[3]), .f(L4[3]), .cout(C4[3]));
    adder_1 adder4_4(.a(X[4] & Y[4]), .b(L3[5]), .cin(C3[4]), .f(L4[4]), .cout(C4[4]));
    adder_1 adder4_5(.a(X[5] & Y[4]), .b(L3[6]), .cin(C3[5]), .f(L4[5]), .cout(C4[5]));
    adder_1 adder4_6(.a(X[6] & Y[4]), .b(L3[7]), .cin(C3[6]), .f(L4[6]), .cout(C4[6]));
    adder_1 adder4_7(.a(X[7] & Y[4]), .b(L3[8]), .cin(C3[7]), .f(L4[7]), .cout(C4[7]));
    adder_1 adder4_8(.a(X[8] & Y[4]), .b(L3[9]), .cin(C3[8]), .f(L4[8]), .cout(C4[8]));
    adder_1 adder4_9(.a(X[9] & Y[4]), .b(L3[10]), .cin(C3[9]), .f(L4[9]), .cout(C4[9]));
    adder_1 adder4_10(.a(X[10] & Y[4]), .b(L3[11]), .cin(C3[10]), .f(L4[10]), .cout(C4[10]));
    adder_1 adder4_11(.a(X[11] & Y[4]), .b(L3[12]), .cin(C3[11]), .f(L4[11]), .cout(C4[11]));
    adder_1 adder4_12(.a(X[12] & Y[4]), .b(L3[13]), .cin(C3[12]), .f(L4[12]), .cout(C4[12]));
    adder_1 adder4_13(.a(X[13] & Y[4]), .b(L3[14]), .cin(C3[13]), .f(L4[13]), .cout(C4[13]));
    adder_1 adder4_14(.a(X[14] & Y[4]), .b(L3[15]), .cin(C3[14]), .f(L4[14]), .cout(C4[14]));
    adder_1 adder4_15(.a(X[15] & Y[4]), .b(L3[16]), .cin(C3[15]), .f(L4[15]), .cout(C4[15]));
    adder_1 adder4_16(.a(X[16] & Y[4]), .b(L3[17]), .cin(C3[16]), .f(L4[16]), .cout(C4[16]));
    adder_1 adder4_17(.a(X[17] & Y[4]), .b(L3[18]), .cin(C3[17]), .f(L4[17]), .cout(C4[17]));
    adder_1 adder4_18(.a(X[18] & Y[4]), .b(L3[19]), .cin(C3[18]), .f(L4[18]), .cout(C4[18]));
    adder_1 adder4_19(.a(X[19] & Y[4]), .b(L3[20]), .cin(C3[19]), .f(L4[19]), .cout(C4[19]));
    adder_1 adder4_20(.a(X[20] & Y[4]), .b(L3[21]), .cin(C3[20]), .f(L4[20]), .cout(C4[20]));
    adder_1 adder4_21(.a(X[21] & Y[4]), .b(L3[22]), .cin(C3[21]), .f(L4[21]), .cout(C4[21]));
    adder_1 adder4_22(.a(X[22] & Y[4]), .b(L3[23]), .cin(C3[22]), .f(L4[22]), .cout(C4[22]));
    adder_1 adder4_23(.a(X[23] & Y[4]), .b(L3[24]), .cin(C3[23]), .f(L4[23]), .cout(C4[23]));
    adder_1 adder4_24(.a(X[24] & Y[4]), .b(L3[25]), .cin(C3[24]), .f(L4[24]), .cout(C4[24]));
    adder_1 adder4_25(.a(X[25] & Y[4]), .b(L3[26]), .cin(C3[25]), .f(L4[25]), .cout(C4[25]));
    adder_1 adder4_26(.a(X[26] & Y[4]), .b(L3[27]), .cin(C3[26]), .f(L4[26]), .cout(C4[26]));
    adder_1 adder4_27(.a(X[27] & Y[4]), .b(L3[28]), .cin(C3[27]), .f(L4[27]), .cout(C4[27]));
    adder_1 adder4_28(.a(X[28] & Y[4]), .b(L3[29]), .cin(C3[28]), .f(L4[28]), .cout(C4[28]));
    adder_1 adder4_29(.a(X[29] & Y[4]), .b(L3[30]), .cin(C3[29]), .f(L4[29]), .cout(C4[29]));
    adder_1 adder4_30(.a(X[30] & Y[4]), .b(L3[31]), .cin(C3[30]), .f(L4[30]), .cout(C4[30]));
    assign L4[31] = X[31] & Y[4];
    wire [31:0] L5, C5;
    adder_1 adder5_0(.a(X[0] & Y[5]), .b(L4[1]), .cin(C4[0]), .f(L5[0]), .cout(C5[0]));
    adder_1 adder5_1(.a(X[1] & Y[5]), .b(L4[2]), .cin(C4[1]), .f(L5[1]), .cout(C5[1]));
    adder_1 adder5_2(.a(X[2] & Y[5]), .b(L4[3]), .cin(C4[2]), .f(L5[2]), .cout(C5[2]));
    adder_1 adder5_3(.a(X[3] & Y[5]), .b(L4[4]), .cin(C4[3]), .f(L5[3]), .cout(C5[3]));
    adder_1 adder5_4(.a(X[4] & Y[5]), .b(L4[5]), .cin(C4[4]), .f(L5[4]), .cout(C5[4]));
    adder_1 adder5_5(.a(X[5] & Y[5]), .b(L4[6]), .cin(C4[5]), .f(L5[5]), .cout(C5[5]));
    adder_1 adder5_6(.a(X[6] & Y[5]), .b(L4[7]), .cin(C4[6]), .f(L5[6]), .cout(C5[6]));
    adder_1 adder5_7(.a(X[7] & Y[5]), .b(L4[8]), .cin(C4[7]), .f(L5[7]), .cout(C5[7]));
    adder_1 adder5_8(.a(X[8] & Y[5]), .b(L4[9]), .cin(C4[8]), .f(L5[8]), .cout(C5[8]));
    adder_1 adder5_9(.a(X[9] & Y[5]), .b(L4[10]), .cin(C4[9]), .f(L5[9]), .cout(C5[9]));
    adder_1 adder5_10(.a(X[10] & Y[5]), .b(L4[11]), .cin(C4[10]), .f(L5[10]), .cout(C5[10]));
    adder_1 adder5_11(.a(X[11] & Y[5]), .b(L4[12]), .cin(C4[11]), .f(L5[11]), .cout(C5[11]));
    adder_1 adder5_12(.a(X[12] & Y[5]), .b(L4[13]), .cin(C4[12]), .f(L5[12]), .cout(C5[12]));
    adder_1 adder5_13(.a(X[13] & Y[5]), .b(L4[14]), .cin(C4[13]), .f(L5[13]), .cout(C5[13]));
    adder_1 adder5_14(.a(X[14] & Y[5]), .b(L4[15]), .cin(C4[14]), .f(L5[14]), .cout(C5[14]));
    adder_1 adder5_15(.a(X[15] & Y[5]), .b(L4[16]), .cin(C4[15]), .f(L5[15]), .cout(C5[15]));
    adder_1 adder5_16(.a(X[16] & Y[5]), .b(L4[17]), .cin(C4[16]), .f(L5[16]), .cout(C5[16]));
    adder_1 adder5_17(.a(X[17] & Y[5]), .b(L4[18]), .cin(C4[17]), .f(L5[17]), .cout(C5[17]));
    adder_1 adder5_18(.a(X[18] & Y[5]), .b(L4[19]), .cin(C4[18]), .f(L5[18]), .cout(C5[18]));
    adder_1 adder5_19(.a(X[19] & Y[5]), .b(L4[20]), .cin(C4[19]), .f(L5[19]), .cout(C5[19]));
    adder_1 adder5_20(.a(X[20] & Y[5]), .b(L4[21]), .cin(C4[20]), .f(L5[20]), .cout(C5[20]));
    adder_1 adder5_21(.a(X[21] & Y[5]), .b(L4[22]), .cin(C4[21]), .f(L5[21]), .cout(C5[21]));
    adder_1 adder5_22(.a(X[22] & Y[5]), .b(L4[23]), .cin(C4[22]), .f(L5[22]), .cout(C5[22]));
    adder_1 adder5_23(.a(X[23] & Y[5]), .b(L4[24]), .cin(C4[23]), .f(L5[23]), .cout(C5[23]));
    adder_1 adder5_24(.a(X[24] & Y[5]), .b(L4[25]), .cin(C4[24]), .f(L5[24]), .cout(C5[24]));
    adder_1 adder5_25(.a(X[25] & Y[5]), .b(L4[26]), .cin(C4[25]), .f(L5[25]), .cout(C5[25]));
    adder_1 adder5_26(.a(X[26] & Y[5]), .b(L4[27]), .cin(C4[26]), .f(L5[26]), .cout(C5[26]));
    adder_1 adder5_27(.a(X[27] & Y[5]), .b(L4[28]), .cin(C4[27]), .f(L5[27]), .cout(C5[27]));
    adder_1 adder5_28(.a(X[28] & Y[5]), .b(L4[29]), .cin(C4[28]), .f(L5[28]), .cout(C5[28]));
    adder_1 adder5_29(.a(X[29] & Y[5]), .b(L4[30]), .cin(C4[29]), .f(L5[29]), .cout(C5[29]));
    adder_1 adder5_30(.a(X[30] & Y[5]), .b(L4[31]), .cin(C4[30]), .f(L5[30]), .cout(C5[30]));
    assign L5[31] = X[31] & Y[5];
    wire [31:0] L6, C6;
    adder_1 adder6_0(.a(X[0] & Y[6]), .b(L5[1]), .cin(C5[0]), .f(L6[0]), .cout(C6[0]));
    adder_1 adder6_1(.a(X[1] & Y[6]), .b(L5[2]), .cin(C5[1]), .f(L6[1]), .cout(C6[1]));
    adder_1 adder6_2(.a(X[2] & Y[6]), .b(L5[3]), .cin(C5[2]), .f(L6[2]), .cout(C6[2]));
    adder_1 adder6_3(.a(X[3] & Y[6]), .b(L5[4]), .cin(C5[3]), .f(L6[3]), .cout(C6[3]));
    adder_1 adder6_4(.a(X[4] & Y[6]), .b(L5[5]), .cin(C5[4]), .f(L6[4]), .cout(C6[4]));
    adder_1 adder6_5(.a(X[5] & Y[6]), .b(L5[6]), .cin(C5[5]), .f(L6[5]), .cout(C6[5]));
    adder_1 adder6_6(.a(X[6] & Y[6]), .b(L5[7]), .cin(C5[6]), .f(L6[6]), .cout(C6[6]));
    adder_1 adder6_7(.a(X[7] & Y[6]), .b(L5[8]), .cin(C5[7]), .f(L6[7]), .cout(C6[7]));
    adder_1 adder6_8(.a(X[8] & Y[6]), .b(L5[9]), .cin(C5[8]), .f(L6[8]), .cout(C6[8]));
    adder_1 adder6_9(.a(X[9] & Y[6]), .b(L5[10]), .cin(C5[9]), .f(L6[9]), .cout(C6[9]));
    adder_1 adder6_10(.a(X[10] & Y[6]), .b(L5[11]), .cin(C5[10]), .f(L6[10]), .cout(C6[10]));
    adder_1 adder6_11(.a(X[11] & Y[6]), .b(L5[12]), .cin(C5[11]), .f(L6[11]), .cout(C6[11]));
    adder_1 adder6_12(.a(X[12] & Y[6]), .b(L5[13]), .cin(C5[12]), .f(L6[12]), .cout(C6[12]));
    adder_1 adder6_13(.a(X[13] & Y[6]), .b(L5[14]), .cin(C5[13]), .f(L6[13]), .cout(C6[13]));
    adder_1 adder6_14(.a(X[14] & Y[6]), .b(L5[15]), .cin(C5[14]), .f(L6[14]), .cout(C6[14]));
    adder_1 adder6_15(.a(X[15] & Y[6]), .b(L5[16]), .cin(C5[15]), .f(L6[15]), .cout(C6[15]));
    adder_1 adder6_16(.a(X[16] & Y[6]), .b(L5[17]), .cin(C5[16]), .f(L6[16]), .cout(C6[16]));
    adder_1 adder6_17(.a(X[17] & Y[6]), .b(L5[18]), .cin(C5[17]), .f(L6[17]), .cout(C6[17]));
    adder_1 adder6_18(.a(X[18] & Y[6]), .b(L5[19]), .cin(C5[18]), .f(L6[18]), .cout(C6[18]));
    adder_1 adder6_19(.a(X[19] & Y[6]), .b(L5[20]), .cin(C5[19]), .f(L6[19]), .cout(C6[19]));
    adder_1 adder6_20(.a(X[20] & Y[6]), .b(L5[21]), .cin(C5[20]), .f(L6[20]), .cout(C6[20]));
    adder_1 adder6_21(.a(X[21] & Y[6]), .b(L5[22]), .cin(C5[21]), .f(L6[21]), .cout(C6[21]));
    adder_1 adder6_22(.a(X[22] & Y[6]), .b(L5[23]), .cin(C5[22]), .f(L6[22]), .cout(C6[22]));
    adder_1 adder6_23(.a(X[23] & Y[6]), .b(L5[24]), .cin(C5[23]), .f(L6[23]), .cout(C6[23]));
    adder_1 adder6_24(.a(X[24] & Y[6]), .b(L5[25]), .cin(C5[24]), .f(L6[24]), .cout(C6[24]));
    adder_1 adder6_25(.a(X[25] & Y[6]), .b(L5[26]), .cin(C5[25]), .f(L6[25]), .cout(C6[25]));
    adder_1 adder6_26(.a(X[26] & Y[6]), .b(L5[27]), .cin(C5[26]), .f(L6[26]), .cout(C6[26]));
    adder_1 adder6_27(.a(X[27] & Y[6]), .b(L5[28]), .cin(C5[27]), .f(L6[27]), .cout(C6[27]));
    adder_1 adder6_28(.a(X[28] & Y[6]), .b(L5[29]), .cin(C5[28]), .f(L6[28]), .cout(C6[28]));
    adder_1 adder6_29(.a(X[29] & Y[6]), .b(L5[30]), .cin(C5[29]), .f(L6[29]), .cout(C6[29]));
    adder_1 adder6_30(.a(X[30] & Y[6]), .b(L5[31]), .cin(C5[30]), .f(L6[30]), .cout(C6[30]));
    assign L6[31] = X[31] & Y[6];
    wire [31:0] L7, C7;
    adder_1 adder7_0(.a(X[0] & Y[7]), .b(L6[1]), .cin(C6[0]), .f(L7[0]), .cout(C7[0]));
    adder_1 adder7_1(.a(X[1] & Y[7]), .b(L6[2]), .cin(C6[1]), .f(L7[1]), .cout(C7[1]));
    adder_1 adder7_2(.a(X[2] & Y[7]), .b(L6[3]), .cin(C6[2]), .f(L7[2]), .cout(C7[2]));
    adder_1 adder7_3(.a(X[3] & Y[7]), .b(L6[4]), .cin(C6[3]), .f(L7[3]), .cout(C7[3]));
    adder_1 adder7_4(.a(X[4] & Y[7]), .b(L6[5]), .cin(C6[4]), .f(L7[4]), .cout(C7[4]));
    adder_1 adder7_5(.a(X[5] & Y[7]), .b(L6[6]), .cin(C6[5]), .f(L7[5]), .cout(C7[5]));
    adder_1 adder7_6(.a(X[6] & Y[7]), .b(L6[7]), .cin(C6[6]), .f(L7[6]), .cout(C7[6]));
    adder_1 adder7_7(.a(X[7] & Y[7]), .b(L6[8]), .cin(C6[7]), .f(L7[7]), .cout(C7[7]));
    adder_1 adder7_8(.a(X[8] & Y[7]), .b(L6[9]), .cin(C6[8]), .f(L7[8]), .cout(C7[8]));
    adder_1 adder7_9(.a(X[9] & Y[7]), .b(L6[10]), .cin(C6[9]), .f(L7[9]), .cout(C7[9]));
    adder_1 adder7_10(.a(X[10] & Y[7]), .b(L6[11]), .cin(C6[10]), .f(L7[10]), .cout(C7[10]));
    adder_1 adder7_11(.a(X[11] & Y[7]), .b(L6[12]), .cin(C6[11]), .f(L7[11]), .cout(C7[11]));
    adder_1 adder7_12(.a(X[12] & Y[7]), .b(L6[13]), .cin(C6[12]), .f(L7[12]), .cout(C7[12]));
    adder_1 adder7_13(.a(X[13] & Y[7]), .b(L6[14]), .cin(C6[13]), .f(L7[13]), .cout(C7[13]));
    adder_1 adder7_14(.a(X[14] & Y[7]), .b(L6[15]), .cin(C6[14]), .f(L7[14]), .cout(C7[14]));
    adder_1 adder7_15(.a(X[15] & Y[7]), .b(L6[16]), .cin(C6[15]), .f(L7[15]), .cout(C7[15]));
    adder_1 adder7_16(.a(X[16] & Y[7]), .b(L6[17]), .cin(C6[16]), .f(L7[16]), .cout(C7[16]));
    adder_1 adder7_17(.a(X[17] & Y[7]), .b(L6[18]), .cin(C6[17]), .f(L7[17]), .cout(C7[17]));
    adder_1 adder7_18(.a(X[18] & Y[7]), .b(L6[19]), .cin(C6[18]), .f(L7[18]), .cout(C7[18]));
    adder_1 adder7_19(.a(X[19] & Y[7]), .b(L6[20]), .cin(C6[19]), .f(L7[19]), .cout(C7[19]));
    adder_1 adder7_20(.a(X[20] & Y[7]), .b(L6[21]), .cin(C6[20]), .f(L7[20]), .cout(C7[20]));
    adder_1 adder7_21(.a(X[21] & Y[7]), .b(L6[22]), .cin(C6[21]), .f(L7[21]), .cout(C7[21]));
    adder_1 adder7_22(.a(X[22] & Y[7]), .b(L6[23]), .cin(C6[22]), .f(L7[22]), .cout(C7[22]));
    adder_1 adder7_23(.a(X[23] & Y[7]), .b(L6[24]), .cin(C6[23]), .f(L7[23]), .cout(C7[23]));
    adder_1 adder7_24(.a(X[24] & Y[7]), .b(L6[25]), .cin(C6[24]), .f(L7[24]), .cout(C7[24]));
    adder_1 adder7_25(.a(X[25] & Y[7]), .b(L6[26]), .cin(C6[25]), .f(L7[25]), .cout(C7[25]));
    adder_1 adder7_26(.a(X[26] & Y[7]), .b(L6[27]), .cin(C6[26]), .f(L7[26]), .cout(C7[26]));
    adder_1 adder7_27(.a(X[27] & Y[7]), .b(L6[28]), .cin(C6[27]), .f(L7[27]), .cout(C7[27]));
    adder_1 adder7_28(.a(X[28] & Y[7]), .b(L6[29]), .cin(C6[28]), .f(L7[28]), .cout(C7[28]));
    adder_1 adder7_29(.a(X[29] & Y[7]), .b(L6[30]), .cin(C6[29]), .f(L7[29]), .cout(C7[29]));
    adder_1 adder7_30(.a(X[30] & Y[7]), .b(L6[31]), .cin(C6[30]), .f(L7[30]), .cout(C7[30]));
    assign L7[31] = X[31] & Y[7];
    wire [31:0] L8, C8;
    adder_1 adder8_0(.a(X[0] & Y[8]), .b(L7[1]), .cin(C7[0]), .f(L8[0]), .cout(C8[0]));
    adder_1 adder8_1(.a(X[1] & Y[8]), .b(L7[2]), .cin(C7[1]), .f(L8[1]), .cout(C8[1]));
    adder_1 adder8_2(.a(X[2] & Y[8]), .b(L7[3]), .cin(C7[2]), .f(L8[2]), .cout(C8[2]));
    adder_1 adder8_3(.a(X[3] & Y[8]), .b(L7[4]), .cin(C7[3]), .f(L8[3]), .cout(C8[3]));
    adder_1 adder8_4(.a(X[4] & Y[8]), .b(L7[5]), .cin(C7[4]), .f(L8[4]), .cout(C8[4]));
    adder_1 adder8_5(.a(X[5] & Y[8]), .b(L7[6]), .cin(C7[5]), .f(L8[5]), .cout(C8[5]));
    adder_1 adder8_6(.a(X[6] & Y[8]), .b(L7[7]), .cin(C7[6]), .f(L8[6]), .cout(C8[6]));
    adder_1 adder8_7(.a(X[7] & Y[8]), .b(L7[8]), .cin(C7[7]), .f(L8[7]), .cout(C8[7]));
    adder_1 adder8_8(.a(X[8] & Y[8]), .b(L7[9]), .cin(C7[8]), .f(L8[8]), .cout(C8[8]));
    adder_1 adder8_9(.a(X[9] & Y[8]), .b(L7[10]), .cin(C7[9]), .f(L8[9]), .cout(C8[9]));
    adder_1 adder8_10(.a(X[10] & Y[8]), .b(L7[11]), .cin(C7[10]), .f(L8[10]), .cout(C8[10]));
    adder_1 adder8_11(.a(X[11] & Y[8]), .b(L7[12]), .cin(C7[11]), .f(L8[11]), .cout(C8[11]));
    adder_1 adder8_12(.a(X[12] & Y[8]), .b(L7[13]), .cin(C7[12]), .f(L8[12]), .cout(C8[12]));
    adder_1 adder8_13(.a(X[13] & Y[8]), .b(L7[14]), .cin(C7[13]), .f(L8[13]), .cout(C8[13]));
    adder_1 adder8_14(.a(X[14] & Y[8]), .b(L7[15]), .cin(C7[14]), .f(L8[14]), .cout(C8[14]));
    adder_1 adder8_15(.a(X[15] & Y[8]), .b(L7[16]), .cin(C7[15]), .f(L8[15]), .cout(C8[15]));
    adder_1 adder8_16(.a(X[16] & Y[8]), .b(L7[17]), .cin(C7[16]), .f(L8[16]), .cout(C8[16]));
    adder_1 adder8_17(.a(X[17] & Y[8]), .b(L7[18]), .cin(C7[17]), .f(L8[17]), .cout(C8[17]));
    adder_1 adder8_18(.a(X[18] & Y[8]), .b(L7[19]), .cin(C7[18]), .f(L8[18]), .cout(C8[18]));
    adder_1 adder8_19(.a(X[19] & Y[8]), .b(L7[20]), .cin(C7[19]), .f(L8[19]), .cout(C8[19]));
    adder_1 adder8_20(.a(X[20] & Y[8]), .b(L7[21]), .cin(C7[20]), .f(L8[20]), .cout(C8[20]));
    adder_1 adder8_21(.a(X[21] & Y[8]), .b(L7[22]), .cin(C7[21]), .f(L8[21]), .cout(C8[21]));
    adder_1 adder8_22(.a(X[22] & Y[8]), .b(L7[23]), .cin(C7[22]), .f(L8[22]), .cout(C8[22]));
    adder_1 adder8_23(.a(X[23] & Y[8]), .b(L7[24]), .cin(C7[23]), .f(L8[23]), .cout(C8[23]));
    adder_1 adder8_24(.a(X[24] & Y[8]), .b(L7[25]), .cin(C7[24]), .f(L8[24]), .cout(C8[24]));
    adder_1 adder8_25(.a(X[25] & Y[8]), .b(L7[26]), .cin(C7[25]), .f(L8[25]), .cout(C8[25]));
    adder_1 adder8_26(.a(X[26] & Y[8]), .b(L7[27]), .cin(C7[26]), .f(L8[26]), .cout(C8[26]));
    adder_1 adder8_27(.a(X[27] & Y[8]), .b(L7[28]), .cin(C7[27]), .f(L8[27]), .cout(C8[27]));
    adder_1 adder8_28(.a(X[28] & Y[8]), .b(L7[29]), .cin(C7[28]), .f(L8[28]), .cout(C8[28]));
    adder_1 adder8_29(.a(X[29] & Y[8]), .b(L7[30]), .cin(C7[29]), .f(L8[29]), .cout(C8[29]));
    adder_1 adder8_30(.a(X[30] & Y[8]), .b(L7[31]), .cin(C7[30]), .f(L8[30]), .cout(C8[30]));
    assign L8[31] = X[31] & Y[8];
    wire [31:0] L9, C9;
    adder_1 adder9_0(.a(X[0] & Y[9]), .b(L8[1]), .cin(C8[0]), .f(L9[0]), .cout(C9[0]));
    adder_1 adder9_1(.a(X[1] & Y[9]), .b(L8[2]), .cin(C8[1]), .f(L9[1]), .cout(C9[1]));
    adder_1 adder9_2(.a(X[2] & Y[9]), .b(L8[3]), .cin(C8[2]), .f(L9[2]), .cout(C9[2]));
    adder_1 adder9_3(.a(X[3] & Y[9]), .b(L8[4]), .cin(C8[3]), .f(L9[3]), .cout(C9[3]));
    adder_1 adder9_4(.a(X[4] & Y[9]), .b(L8[5]), .cin(C8[4]), .f(L9[4]), .cout(C9[4]));
    adder_1 adder9_5(.a(X[5] & Y[9]), .b(L8[6]), .cin(C8[5]), .f(L9[5]), .cout(C9[5]));
    adder_1 adder9_6(.a(X[6] & Y[9]), .b(L8[7]), .cin(C8[6]), .f(L9[6]), .cout(C9[6]));
    adder_1 adder9_7(.a(X[7] & Y[9]), .b(L8[8]), .cin(C8[7]), .f(L9[7]), .cout(C9[7]));
    adder_1 adder9_8(.a(X[8] & Y[9]), .b(L8[9]), .cin(C8[8]), .f(L9[8]), .cout(C9[8]));
    adder_1 adder9_9(.a(X[9] & Y[9]), .b(L8[10]), .cin(C8[9]), .f(L9[9]), .cout(C9[9]));
    adder_1 adder9_10(.a(X[10] & Y[9]), .b(L8[11]), .cin(C8[10]), .f(L9[10]), .cout(C9[10]));
    adder_1 adder9_11(.a(X[11] & Y[9]), .b(L8[12]), .cin(C8[11]), .f(L9[11]), .cout(C9[11]));
    adder_1 adder9_12(.a(X[12] & Y[9]), .b(L8[13]), .cin(C8[12]), .f(L9[12]), .cout(C9[12]));
    adder_1 adder9_13(.a(X[13] & Y[9]), .b(L8[14]), .cin(C8[13]), .f(L9[13]), .cout(C9[13]));
    adder_1 adder9_14(.a(X[14] & Y[9]), .b(L8[15]), .cin(C8[14]), .f(L9[14]), .cout(C9[14]));
    adder_1 adder9_15(.a(X[15] & Y[9]), .b(L8[16]), .cin(C8[15]), .f(L9[15]), .cout(C9[15]));
    adder_1 adder9_16(.a(X[16] & Y[9]), .b(L8[17]), .cin(C8[16]), .f(L9[16]), .cout(C9[16]));
    adder_1 adder9_17(.a(X[17] & Y[9]), .b(L8[18]), .cin(C8[17]), .f(L9[17]), .cout(C9[17]));
    adder_1 adder9_18(.a(X[18] & Y[9]), .b(L8[19]), .cin(C8[18]), .f(L9[18]), .cout(C9[18]));
    adder_1 adder9_19(.a(X[19] & Y[9]), .b(L8[20]), .cin(C8[19]), .f(L9[19]), .cout(C9[19]));
    adder_1 adder9_20(.a(X[20] & Y[9]), .b(L8[21]), .cin(C8[20]), .f(L9[20]), .cout(C9[20]));
    adder_1 adder9_21(.a(X[21] & Y[9]), .b(L8[22]), .cin(C8[21]), .f(L9[21]), .cout(C9[21]));
    adder_1 adder9_22(.a(X[22] & Y[9]), .b(L8[23]), .cin(C8[22]), .f(L9[22]), .cout(C9[22]));
    adder_1 adder9_23(.a(X[23] & Y[9]), .b(L8[24]), .cin(C8[23]), .f(L9[23]), .cout(C9[23]));
    adder_1 adder9_24(.a(X[24] & Y[9]), .b(L8[25]), .cin(C8[24]), .f(L9[24]), .cout(C9[24]));
    adder_1 adder9_25(.a(X[25] & Y[9]), .b(L8[26]), .cin(C8[25]), .f(L9[25]), .cout(C9[25]));
    adder_1 adder9_26(.a(X[26] & Y[9]), .b(L8[27]), .cin(C8[26]), .f(L9[26]), .cout(C9[26]));
    adder_1 adder9_27(.a(X[27] & Y[9]), .b(L8[28]), .cin(C8[27]), .f(L9[27]), .cout(C9[27]));
    adder_1 adder9_28(.a(X[28] & Y[9]), .b(L8[29]), .cin(C8[28]), .f(L9[28]), .cout(C9[28]));
    adder_1 adder9_29(.a(X[29] & Y[9]), .b(L8[30]), .cin(C8[29]), .f(L9[29]), .cout(C9[29]));
    adder_1 adder9_30(.a(X[30] & Y[9]), .b(L8[31]), .cin(C8[30]), .f(L9[30]), .cout(C9[30]));
    assign L9[31] = X[31] & Y[9];
    wire [31:0] L10, C10;
    adder_1 adder10_0(.a(X[0] & Y[10]), .b(L9[1]), .cin(C9[0]), .f(L10[0]), .cout(C10[0]));
    adder_1 adder10_1(.a(X[1] & Y[10]), .b(L9[2]), .cin(C9[1]), .f(L10[1]), .cout(C10[1]));
    adder_1 adder10_2(.a(X[2] & Y[10]), .b(L9[3]), .cin(C9[2]), .f(L10[2]), .cout(C10[2]));
    adder_1 adder10_3(.a(X[3] & Y[10]), .b(L9[4]), .cin(C9[3]), .f(L10[3]), .cout(C10[3]));
    adder_1 adder10_4(.a(X[4] & Y[10]), .b(L9[5]), .cin(C9[4]), .f(L10[4]), .cout(C10[4]));
    adder_1 adder10_5(.a(X[5] & Y[10]), .b(L9[6]), .cin(C9[5]), .f(L10[5]), .cout(C10[5]));
    adder_1 adder10_6(.a(X[6] & Y[10]), .b(L9[7]), .cin(C9[6]), .f(L10[6]), .cout(C10[6]));
    adder_1 adder10_7(.a(X[7] & Y[10]), .b(L9[8]), .cin(C9[7]), .f(L10[7]), .cout(C10[7]));
    adder_1 adder10_8(.a(X[8] & Y[10]), .b(L9[9]), .cin(C9[8]), .f(L10[8]), .cout(C10[8]));
    adder_1 adder10_9(.a(X[9] & Y[10]), .b(L9[10]), .cin(C9[9]), .f(L10[9]), .cout(C10[9]));
    adder_1 adder10_10(.a(X[10] & Y[10]), .b(L9[11]), .cin(C9[10]), .f(L10[10]), .cout(C10[10]));
    adder_1 adder10_11(.a(X[11] & Y[10]), .b(L9[12]), .cin(C9[11]), .f(L10[11]), .cout(C10[11]));
    adder_1 adder10_12(.a(X[12] & Y[10]), .b(L9[13]), .cin(C9[12]), .f(L10[12]), .cout(C10[12]));
    adder_1 adder10_13(.a(X[13] & Y[10]), .b(L9[14]), .cin(C9[13]), .f(L10[13]), .cout(C10[13]));
    adder_1 adder10_14(.a(X[14] & Y[10]), .b(L9[15]), .cin(C9[14]), .f(L10[14]), .cout(C10[14]));
    adder_1 adder10_15(.a(X[15] & Y[10]), .b(L9[16]), .cin(C9[15]), .f(L10[15]), .cout(C10[15]));
    adder_1 adder10_16(.a(X[16] & Y[10]), .b(L9[17]), .cin(C9[16]), .f(L10[16]), .cout(C10[16]));
    adder_1 adder10_17(.a(X[17] & Y[10]), .b(L9[18]), .cin(C9[17]), .f(L10[17]), .cout(C10[17]));
    adder_1 adder10_18(.a(X[18] & Y[10]), .b(L9[19]), .cin(C9[18]), .f(L10[18]), .cout(C10[18]));
    adder_1 adder10_19(.a(X[19] & Y[10]), .b(L9[20]), .cin(C9[19]), .f(L10[19]), .cout(C10[19]));
    adder_1 adder10_20(.a(X[20] & Y[10]), .b(L9[21]), .cin(C9[20]), .f(L10[20]), .cout(C10[20]));
    adder_1 adder10_21(.a(X[21] & Y[10]), .b(L9[22]), .cin(C9[21]), .f(L10[21]), .cout(C10[21]));
    adder_1 adder10_22(.a(X[22] & Y[10]), .b(L9[23]), .cin(C9[22]), .f(L10[22]), .cout(C10[22]));
    adder_1 adder10_23(.a(X[23] & Y[10]), .b(L9[24]), .cin(C9[23]), .f(L10[23]), .cout(C10[23]));
    adder_1 adder10_24(.a(X[24] & Y[10]), .b(L9[25]), .cin(C9[24]), .f(L10[24]), .cout(C10[24]));
    adder_1 adder10_25(.a(X[25] & Y[10]), .b(L9[26]), .cin(C9[25]), .f(L10[25]), .cout(C10[25]));
    adder_1 adder10_26(.a(X[26] & Y[10]), .b(L9[27]), .cin(C9[26]), .f(L10[26]), .cout(C10[26]));
    adder_1 adder10_27(.a(X[27] & Y[10]), .b(L9[28]), .cin(C9[27]), .f(L10[27]), .cout(C10[27]));
    adder_1 adder10_28(.a(X[28] & Y[10]), .b(L9[29]), .cin(C9[28]), .f(L10[28]), .cout(C10[28]));
    adder_1 adder10_29(.a(X[29] & Y[10]), .b(L9[30]), .cin(C9[29]), .f(L10[29]), .cout(C10[29]));
    adder_1 adder10_30(.a(X[30] & Y[10]), .b(L9[31]), .cin(C9[30]), .f(L10[30]), .cout(C10[30]));
    assign L10[31] = X[31] & Y[10];
    wire [31:0] L11, C11;
    adder_1 adder11_0(.a(X[0] & Y[11]), .b(L10[1]), .cin(C10[0]), .f(L11[0]), .cout(C11[0]));
    adder_1 adder11_1(.a(X[1] & Y[11]), .b(L10[2]), .cin(C10[1]), .f(L11[1]), .cout(C11[1]));
    adder_1 adder11_2(.a(X[2] & Y[11]), .b(L10[3]), .cin(C10[2]), .f(L11[2]), .cout(C11[2]));
    adder_1 adder11_3(.a(X[3] & Y[11]), .b(L10[4]), .cin(C10[3]), .f(L11[3]), .cout(C11[3]));
    adder_1 adder11_4(.a(X[4] & Y[11]), .b(L10[5]), .cin(C10[4]), .f(L11[4]), .cout(C11[4]));
    adder_1 adder11_5(.a(X[5] & Y[11]), .b(L10[6]), .cin(C10[5]), .f(L11[5]), .cout(C11[5]));
    adder_1 adder11_6(.a(X[6] & Y[11]), .b(L10[7]), .cin(C10[6]), .f(L11[6]), .cout(C11[6]));
    adder_1 adder11_7(.a(X[7] & Y[11]), .b(L10[8]), .cin(C10[7]), .f(L11[7]), .cout(C11[7]));
    adder_1 adder11_8(.a(X[8] & Y[11]), .b(L10[9]), .cin(C10[8]), .f(L11[8]), .cout(C11[8]));
    adder_1 adder11_9(.a(X[9] & Y[11]), .b(L10[10]), .cin(C10[9]), .f(L11[9]), .cout(C11[9]));
    adder_1 adder11_10(.a(X[10] & Y[11]), .b(L10[11]), .cin(C10[10]), .f(L11[10]), .cout(C11[10]));
    adder_1 adder11_11(.a(X[11] & Y[11]), .b(L10[12]), .cin(C10[11]), .f(L11[11]), .cout(C11[11]));
    adder_1 adder11_12(.a(X[12] & Y[11]), .b(L10[13]), .cin(C10[12]), .f(L11[12]), .cout(C11[12]));
    adder_1 adder11_13(.a(X[13] & Y[11]), .b(L10[14]), .cin(C10[13]), .f(L11[13]), .cout(C11[13]));
    adder_1 adder11_14(.a(X[14] & Y[11]), .b(L10[15]), .cin(C10[14]), .f(L11[14]), .cout(C11[14]));
    adder_1 adder11_15(.a(X[15] & Y[11]), .b(L10[16]), .cin(C10[15]), .f(L11[15]), .cout(C11[15]));
    adder_1 adder11_16(.a(X[16] & Y[11]), .b(L10[17]), .cin(C10[16]), .f(L11[16]), .cout(C11[16]));
    adder_1 adder11_17(.a(X[17] & Y[11]), .b(L10[18]), .cin(C10[17]), .f(L11[17]), .cout(C11[17]));
    adder_1 adder11_18(.a(X[18] & Y[11]), .b(L10[19]), .cin(C10[18]), .f(L11[18]), .cout(C11[18]));
    adder_1 adder11_19(.a(X[19] & Y[11]), .b(L10[20]), .cin(C10[19]), .f(L11[19]), .cout(C11[19]));
    adder_1 adder11_20(.a(X[20] & Y[11]), .b(L10[21]), .cin(C10[20]), .f(L11[20]), .cout(C11[20]));
    adder_1 adder11_21(.a(X[21] & Y[11]), .b(L10[22]), .cin(C10[21]), .f(L11[21]), .cout(C11[21]));
    adder_1 adder11_22(.a(X[22] & Y[11]), .b(L10[23]), .cin(C10[22]), .f(L11[22]), .cout(C11[22]));
    adder_1 adder11_23(.a(X[23] & Y[11]), .b(L10[24]), .cin(C10[23]), .f(L11[23]), .cout(C11[23]));
    adder_1 adder11_24(.a(X[24] & Y[11]), .b(L10[25]), .cin(C10[24]), .f(L11[24]), .cout(C11[24]));
    adder_1 adder11_25(.a(X[25] & Y[11]), .b(L10[26]), .cin(C10[25]), .f(L11[25]), .cout(C11[25]));
    adder_1 adder11_26(.a(X[26] & Y[11]), .b(L10[27]), .cin(C10[26]), .f(L11[26]), .cout(C11[26]));
    adder_1 adder11_27(.a(X[27] & Y[11]), .b(L10[28]), .cin(C10[27]), .f(L11[27]), .cout(C11[27]));
    adder_1 adder11_28(.a(X[28] & Y[11]), .b(L10[29]), .cin(C10[28]), .f(L11[28]), .cout(C11[28]));
    adder_1 adder11_29(.a(X[29] & Y[11]), .b(L10[30]), .cin(C10[29]), .f(L11[29]), .cout(C11[29]));
    adder_1 adder11_30(.a(X[30] & Y[11]), .b(L10[31]), .cin(C10[30]), .f(L11[30]), .cout(C11[30]));
    assign L11[31] = X[31] & Y[11];
    wire [31:0] L12, C12;
    adder_1 adder12_0(.a(X[0] & Y[12]), .b(L11[1]), .cin(C11[0]), .f(L12[0]), .cout(C12[0]));
    adder_1 adder12_1(.a(X[1] & Y[12]), .b(L11[2]), .cin(C11[1]), .f(L12[1]), .cout(C12[1]));
    adder_1 adder12_2(.a(X[2] & Y[12]), .b(L11[3]), .cin(C11[2]), .f(L12[2]), .cout(C12[2]));
    adder_1 adder12_3(.a(X[3] & Y[12]), .b(L11[4]), .cin(C11[3]), .f(L12[3]), .cout(C12[3]));
    adder_1 adder12_4(.a(X[4] & Y[12]), .b(L11[5]), .cin(C11[4]), .f(L12[4]), .cout(C12[4]));
    adder_1 adder12_5(.a(X[5] & Y[12]), .b(L11[6]), .cin(C11[5]), .f(L12[5]), .cout(C12[5]));
    adder_1 adder12_6(.a(X[6] & Y[12]), .b(L11[7]), .cin(C11[6]), .f(L12[6]), .cout(C12[6]));
    adder_1 adder12_7(.a(X[7] & Y[12]), .b(L11[8]), .cin(C11[7]), .f(L12[7]), .cout(C12[7]));
    adder_1 adder12_8(.a(X[8] & Y[12]), .b(L11[9]), .cin(C11[8]), .f(L12[8]), .cout(C12[8]));
    adder_1 adder12_9(.a(X[9] & Y[12]), .b(L11[10]), .cin(C11[9]), .f(L12[9]), .cout(C12[9]));
    adder_1 adder12_10(.a(X[10] & Y[12]), .b(L11[11]), .cin(C11[10]), .f(L12[10]), .cout(C12[10]));
    adder_1 adder12_11(.a(X[11] & Y[12]), .b(L11[12]), .cin(C11[11]), .f(L12[11]), .cout(C12[11]));
    adder_1 adder12_12(.a(X[12] & Y[12]), .b(L11[13]), .cin(C11[12]), .f(L12[12]), .cout(C12[12]));
    adder_1 adder12_13(.a(X[13] & Y[12]), .b(L11[14]), .cin(C11[13]), .f(L12[13]), .cout(C12[13]));
    adder_1 adder12_14(.a(X[14] & Y[12]), .b(L11[15]), .cin(C11[14]), .f(L12[14]), .cout(C12[14]));
    adder_1 adder12_15(.a(X[15] & Y[12]), .b(L11[16]), .cin(C11[15]), .f(L12[15]), .cout(C12[15]));
    adder_1 adder12_16(.a(X[16] & Y[12]), .b(L11[17]), .cin(C11[16]), .f(L12[16]), .cout(C12[16]));
    adder_1 adder12_17(.a(X[17] & Y[12]), .b(L11[18]), .cin(C11[17]), .f(L12[17]), .cout(C12[17]));
    adder_1 adder12_18(.a(X[18] & Y[12]), .b(L11[19]), .cin(C11[18]), .f(L12[18]), .cout(C12[18]));
    adder_1 adder12_19(.a(X[19] & Y[12]), .b(L11[20]), .cin(C11[19]), .f(L12[19]), .cout(C12[19]));
    adder_1 adder12_20(.a(X[20] & Y[12]), .b(L11[21]), .cin(C11[20]), .f(L12[20]), .cout(C12[20]));
    adder_1 adder12_21(.a(X[21] & Y[12]), .b(L11[22]), .cin(C11[21]), .f(L12[21]), .cout(C12[21]));
    adder_1 adder12_22(.a(X[22] & Y[12]), .b(L11[23]), .cin(C11[22]), .f(L12[22]), .cout(C12[22]));
    adder_1 adder12_23(.a(X[23] & Y[12]), .b(L11[24]), .cin(C11[23]), .f(L12[23]), .cout(C12[23]));
    adder_1 adder12_24(.a(X[24] & Y[12]), .b(L11[25]), .cin(C11[24]), .f(L12[24]), .cout(C12[24]));
    adder_1 adder12_25(.a(X[25] & Y[12]), .b(L11[26]), .cin(C11[25]), .f(L12[25]), .cout(C12[25]));
    adder_1 adder12_26(.a(X[26] & Y[12]), .b(L11[27]), .cin(C11[26]), .f(L12[26]), .cout(C12[26]));
    adder_1 adder12_27(.a(X[27] & Y[12]), .b(L11[28]), .cin(C11[27]), .f(L12[27]), .cout(C12[27]));
    adder_1 adder12_28(.a(X[28] & Y[12]), .b(L11[29]), .cin(C11[28]), .f(L12[28]), .cout(C12[28]));
    adder_1 adder12_29(.a(X[29] & Y[12]), .b(L11[30]), .cin(C11[29]), .f(L12[29]), .cout(C12[29]));
    adder_1 adder12_30(.a(X[30] & Y[12]), .b(L11[31]), .cin(C11[30]), .f(L12[30]), .cout(C12[30]));
    assign L12[31] = X[31] & Y[12];
    wire [31:0] L13, C13;
    adder_1 adder13_0(.a(X[0] & Y[13]), .b(L12[1]), .cin(C12[0]), .f(L13[0]), .cout(C13[0]));
    adder_1 adder13_1(.a(X[1] & Y[13]), .b(L12[2]), .cin(C12[1]), .f(L13[1]), .cout(C13[1]));
    adder_1 adder13_2(.a(X[2] & Y[13]), .b(L12[3]), .cin(C12[2]), .f(L13[2]), .cout(C13[2]));
    adder_1 adder13_3(.a(X[3] & Y[13]), .b(L12[4]), .cin(C12[3]), .f(L13[3]), .cout(C13[3]));
    adder_1 adder13_4(.a(X[4] & Y[13]), .b(L12[5]), .cin(C12[4]), .f(L13[4]), .cout(C13[4]));
    adder_1 adder13_5(.a(X[5] & Y[13]), .b(L12[6]), .cin(C12[5]), .f(L13[5]), .cout(C13[5]));
    adder_1 adder13_6(.a(X[6] & Y[13]), .b(L12[7]), .cin(C12[6]), .f(L13[6]), .cout(C13[6]));
    adder_1 adder13_7(.a(X[7] & Y[13]), .b(L12[8]), .cin(C12[7]), .f(L13[7]), .cout(C13[7]));
    adder_1 adder13_8(.a(X[8] & Y[13]), .b(L12[9]), .cin(C12[8]), .f(L13[8]), .cout(C13[8]));
    adder_1 adder13_9(.a(X[9] & Y[13]), .b(L12[10]), .cin(C12[9]), .f(L13[9]), .cout(C13[9]));
    adder_1 adder13_10(.a(X[10] & Y[13]), .b(L12[11]), .cin(C12[10]), .f(L13[10]), .cout(C13[10]));
    adder_1 adder13_11(.a(X[11] & Y[13]), .b(L12[12]), .cin(C12[11]), .f(L13[11]), .cout(C13[11]));
    adder_1 adder13_12(.a(X[12] & Y[13]), .b(L12[13]), .cin(C12[12]), .f(L13[12]), .cout(C13[12]));
    adder_1 adder13_13(.a(X[13] & Y[13]), .b(L12[14]), .cin(C12[13]), .f(L13[13]), .cout(C13[13]));
    adder_1 adder13_14(.a(X[14] & Y[13]), .b(L12[15]), .cin(C12[14]), .f(L13[14]), .cout(C13[14]));
    adder_1 adder13_15(.a(X[15] & Y[13]), .b(L12[16]), .cin(C12[15]), .f(L13[15]), .cout(C13[15]));
    adder_1 adder13_16(.a(X[16] & Y[13]), .b(L12[17]), .cin(C12[16]), .f(L13[16]), .cout(C13[16]));
    adder_1 adder13_17(.a(X[17] & Y[13]), .b(L12[18]), .cin(C12[17]), .f(L13[17]), .cout(C13[17]));
    adder_1 adder13_18(.a(X[18] & Y[13]), .b(L12[19]), .cin(C12[18]), .f(L13[18]), .cout(C13[18]));
    adder_1 adder13_19(.a(X[19] & Y[13]), .b(L12[20]), .cin(C12[19]), .f(L13[19]), .cout(C13[19]));
    adder_1 adder13_20(.a(X[20] & Y[13]), .b(L12[21]), .cin(C12[20]), .f(L13[20]), .cout(C13[20]));
    adder_1 adder13_21(.a(X[21] & Y[13]), .b(L12[22]), .cin(C12[21]), .f(L13[21]), .cout(C13[21]));
    adder_1 adder13_22(.a(X[22] & Y[13]), .b(L12[23]), .cin(C12[22]), .f(L13[22]), .cout(C13[22]));
    adder_1 adder13_23(.a(X[23] & Y[13]), .b(L12[24]), .cin(C12[23]), .f(L13[23]), .cout(C13[23]));
    adder_1 adder13_24(.a(X[24] & Y[13]), .b(L12[25]), .cin(C12[24]), .f(L13[24]), .cout(C13[24]));
    adder_1 adder13_25(.a(X[25] & Y[13]), .b(L12[26]), .cin(C12[25]), .f(L13[25]), .cout(C13[25]));
    adder_1 adder13_26(.a(X[26] & Y[13]), .b(L12[27]), .cin(C12[26]), .f(L13[26]), .cout(C13[26]));
    adder_1 adder13_27(.a(X[27] & Y[13]), .b(L12[28]), .cin(C12[27]), .f(L13[27]), .cout(C13[27]));
    adder_1 adder13_28(.a(X[28] & Y[13]), .b(L12[29]), .cin(C12[28]), .f(L13[28]), .cout(C13[28]));
    adder_1 adder13_29(.a(X[29] & Y[13]), .b(L12[30]), .cin(C12[29]), .f(L13[29]), .cout(C13[29]));
    adder_1 adder13_30(.a(X[30] & Y[13]), .b(L12[31]), .cin(C12[30]), .f(L13[30]), .cout(C13[30]));
    assign L13[31] = X[31] & Y[13];
    wire [31:0] L14, C14;
    adder_1 adder14_0(.a(X[0] & Y[14]), .b(L13[1]), .cin(C13[0]), .f(L14[0]), .cout(C14[0]));
    adder_1 adder14_1(.a(X[1] & Y[14]), .b(L13[2]), .cin(C13[1]), .f(L14[1]), .cout(C14[1]));
    adder_1 adder14_2(.a(X[2] & Y[14]), .b(L13[3]), .cin(C13[2]), .f(L14[2]), .cout(C14[2]));
    adder_1 adder14_3(.a(X[3] & Y[14]), .b(L13[4]), .cin(C13[3]), .f(L14[3]), .cout(C14[3]));
    adder_1 adder14_4(.a(X[4] & Y[14]), .b(L13[5]), .cin(C13[4]), .f(L14[4]), .cout(C14[4]));
    adder_1 adder14_5(.a(X[5] & Y[14]), .b(L13[6]), .cin(C13[5]), .f(L14[5]), .cout(C14[5]));
    adder_1 adder14_6(.a(X[6] & Y[14]), .b(L13[7]), .cin(C13[6]), .f(L14[6]), .cout(C14[6]));
    adder_1 adder14_7(.a(X[7] & Y[14]), .b(L13[8]), .cin(C13[7]), .f(L14[7]), .cout(C14[7]));
    adder_1 adder14_8(.a(X[8] & Y[14]), .b(L13[9]), .cin(C13[8]), .f(L14[8]), .cout(C14[8]));
    adder_1 adder14_9(.a(X[9] & Y[14]), .b(L13[10]), .cin(C13[9]), .f(L14[9]), .cout(C14[9]));
    adder_1 adder14_10(.a(X[10] & Y[14]), .b(L13[11]), .cin(C13[10]), .f(L14[10]), .cout(C14[10]));
    adder_1 adder14_11(.a(X[11] & Y[14]), .b(L13[12]), .cin(C13[11]), .f(L14[11]), .cout(C14[11]));
    adder_1 adder14_12(.a(X[12] & Y[14]), .b(L13[13]), .cin(C13[12]), .f(L14[12]), .cout(C14[12]));
    adder_1 adder14_13(.a(X[13] & Y[14]), .b(L13[14]), .cin(C13[13]), .f(L14[13]), .cout(C14[13]));
    adder_1 adder14_14(.a(X[14] & Y[14]), .b(L13[15]), .cin(C13[14]), .f(L14[14]), .cout(C14[14]));
    adder_1 adder14_15(.a(X[15] & Y[14]), .b(L13[16]), .cin(C13[15]), .f(L14[15]), .cout(C14[15]));
    adder_1 adder14_16(.a(X[16] & Y[14]), .b(L13[17]), .cin(C13[16]), .f(L14[16]), .cout(C14[16]));
    adder_1 adder14_17(.a(X[17] & Y[14]), .b(L13[18]), .cin(C13[17]), .f(L14[17]), .cout(C14[17]));
    adder_1 adder14_18(.a(X[18] & Y[14]), .b(L13[19]), .cin(C13[18]), .f(L14[18]), .cout(C14[18]));
    adder_1 adder14_19(.a(X[19] & Y[14]), .b(L13[20]), .cin(C13[19]), .f(L14[19]), .cout(C14[19]));
    adder_1 adder14_20(.a(X[20] & Y[14]), .b(L13[21]), .cin(C13[20]), .f(L14[20]), .cout(C14[20]));
    adder_1 adder14_21(.a(X[21] & Y[14]), .b(L13[22]), .cin(C13[21]), .f(L14[21]), .cout(C14[21]));
    adder_1 adder14_22(.a(X[22] & Y[14]), .b(L13[23]), .cin(C13[22]), .f(L14[22]), .cout(C14[22]));
    adder_1 adder14_23(.a(X[23] & Y[14]), .b(L13[24]), .cin(C13[23]), .f(L14[23]), .cout(C14[23]));
    adder_1 adder14_24(.a(X[24] & Y[14]), .b(L13[25]), .cin(C13[24]), .f(L14[24]), .cout(C14[24]));
    adder_1 adder14_25(.a(X[25] & Y[14]), .b(L13[26]), .cin(C13[25]), .f(L14[25]), .cout(C14[25]));
    adder_1 adder14_26(.a(X[26] & Y[14]), .b(L13[27]), .cin(C13[26]), .f(L14[26]), .cout(C14[26]));
    adder_1 adder14_27(.a(X[27] & Y[14]), .b(L13[28]), .cin(C13[27]), .f(L14[27]), .cout(C14[27]));
    adder_1 adder14_28(.a(X[28] & Y[14]), .b(L13[29]), .cin(C13[28]), .f(L14[28]), .cout(C14[28]));
    adder_1 adder14_29(.a(X[29] & Y[14]), .b(L13[30]), .cin(C13[29]), .f(L14[29]), .cout(C14[29]));
    adder_1 adder14_30(.a(X[30] & Y[14]), .b(L13[31]), .cin(C13[30]), .f(L14[30]), .cout(C14[30]));
    assign L14[31] = X[31] & Y[14];
    wire [31:0] L15, C15;
    adder_1 adder15_0(.a(X[0] & Y[15]), .b(L14[1]), .cin(C14[0]), .f(L15[0]), .cout(C15[0]));
    adder_1 adder15_1(.a(X[1] & Y[15]), .b(L14[2]), .cin(C14[1]), .f(L15[1]), .cout(C15[1]));
    adder_1 adder15_2(.a(X[2] & Y[15]), .b(L14[3]), .cin(C14[2]), .f(L15[2]), .cout(C15[2]));
    adder_1 adder15_3(.a(X[3] & Y[15]), .b(L14[4]), .cin(C14[3]), .f(L15[3]), .cout(C15[3]));
    adder_1 adder15_4(.a(X[4] & Y[15]), .b(L14[5]), .cin(C14[4]), .f(L15[4]), .cout(C15[4]));
    adder_1 adder15_5(.a(X[5] & Y[15]), .b(L14[6]), .cin(C14[5]), .f(L15[5]), .cout(C15[5]));
    adder_1 adder15_6(.a(X[6] & Y[15]), .b(L14[7]), .cin(C14[6]), .f(L15[6]), .cout(C15[6]));
    adder_1 adder15_7(.a(X[7] & Y[15]), .b(L14[8]), .cin(C14[7]), .f(L15[7]), .cout(C15[7]));
    adder_1 adder15_8(.a(X[8] & Y[15]), .b(L14[9]), .cin(C14[8]), .f(L15[8]), .cout(C15[8]));
    adder_1 adder15_9(.a(X[9] & Y[15]), .b(L14[10]), .cin(C14[9]), .f(L15[9]), .cout(C15[9]));
    adder_1 adder15_10(.a(X[10] & Y[15]), .b(L14[11]), .cin(C14[10]), .f(L15[10]), .cout(C15[10]));
    adder_1 adder15_11(.a(X[11] & Y[15]), .b(L14[12]), .cin(C14[11]), .f(L15[11]), .cout(C15[11]));
    adder_1 adder15_12(.a(X[12] & Y[15]), .b(L14[13]), .cin(C14[12]), .f(L15[12]), .cout(C15[12]));
    adder_1 adder15_13(.a(X[13] & Y[15]), .b(L14[14]), .cin(C14[13]), .f(L15[13]), .cout(C15[13]));
    adder_1 adder15_14(.a(X[14] & Y[15]), .b(L14[15]), .cin(C14[14]), .f(L15[14]), .cout(C15[14]));
    adder_1 adder15_15(.a(X[15] & Y[15]), .b(L14[16]), .cin(C14[15]), .f(L15[15]), .cout(C15[15]));
    adder_1 adder15_16(.a(X[16] & Y[15]), .b(L14[17]), .cin(C14[16]), .f(L15[16]), .cout(C15[16]));
    adder_1 adder15_17(.a(X[17] & Y[15]), .b(L14[18]), .cin(C14[17]), .f(L15[17]), .cout(C15[17]));
    adder_1 adder15_18(.a(X[18] & Y[15]), .b(L14[19]), .cin(C14[18]), .f(L15[18]), .cout(C15[18]));
    adder_1 adder15_19(.a(X[19] & Y[15]), .b(L14[20]), .cin(C14[19]), .f(L15[19]), .cout(C15[19]));
    adder_1 adder15_20(.a(X[20] & Y[15]), .b(L14[21]), .cin(C14[20]), .f(L15[20]), .cout(C15[20]));
    adder_1 adder15_21(.a(X[21] & Y[15]), .b(L14[22]), .cin(C14[21]), .f(L15[21]), .cout(C15[21]));
    adder_1 adder15_22(.a(X[22] & Y[15]), .b(L14[23]), .cin(C14[22]), .f(L15[22]), .cout(C15[22]));
    adder_1 adder15_23(.a(X[23] & Y[15]), .b(L14[24]), .cin(C14[23]), .f(L15[23]), .cout(C15[23]));
    adder_1 adder15_24(.a(X[24] & Y[15]), .b(L14[25]), .cin(C14[24]), .f(L15[24]), .cout(C15[24]));
    adder_1 adder15_25(.a(X[25] & Y[15]), .b(L14[26]), .cin(C14[25]), .f(L15[25]), .cout(C15[25]));
    adder_1 adder15_26(.a(X[26] & Y[15]), .b(L14[27]), .cin(C14[26]), .f(L15[26]), .cout(C15[26]));
    adder_1 adder15_27(.a(X[27] & Y[15]), .b(L14[28]), .cin(C14[27]), .f(L15[27]), .cout(C15[27]));
    adder_1 adder15_28(.a(X[28] & Y[15]), .b(L14[29]), .cin(C14[28]), .f(L15[28]), .cout(C15[28]));
    adder_1 adder15_29(.a(X[29] & Y[15]), .b(L14[30]), .cin(C14[29]), .f(L15[29]), .cout(C15[29]));
    adder_1 adder15_30(.a(X[30] & Y[15]), .b(L14[31]), .cin(C14[30]), .f(L15[30]), .cout(C15[30]));
    assign L15[31] = X[31] & Y[15];
    wire [31:0] L16, C16;
    adder_1 adder16_0(.a(X[0] & Y[16]), .b(L15[1]), .cin(C15[0]), .f(L16[0]), .cout(C16[0]));
    adder_1 adder16_1(.a(X[1] & Y[16]), .b(L15[2]), .cin(C15[1]), .f(L16[1]), .cout(C16[1]));
    adder_1 adder16_2(.a(X[2] & Y[16]), .b(L15[3]), .cin(C15[2]), .f(L16[2]), .cout(C16[2]));
    adder_1 adder16_3(.a(X[3] & Y[16]), .b(L15[4]), .cin(C15[3]), .f(L16[3]), .cout(C16[3]));
    adder_1 adder16_4(.a(X[4] & Y[16]), .b(L15[5]), .cin(C15[4]), .f(L16[4]), .cout(C16[4]));
    adder_1 adder16_5(.a(X[5] & Y[16]), .b(L15[6]), .cin(C15[5]), .f(L16[5]), .cout(C16[5]));
    adder_1 adder16_6(.a(X[6] & Y[16]), .b(L15[7]), .cin(C15[6]), .f(L16[6]), .cout(C16[6]));
    adder_1 adder16_7(.a(X[7] & Y[16]), .b(L15[8]), .cin(C15[7]), .f(L16[7]), .cout(C16[7]));
    adder_1 adder16_8(.a(X[8] & Y[16]), .b(L15[9]), .cin(C15[8]), .f(L16[8]), .cout(C16[8]));
    adder_1 adder16_9(.a(X[9] & Y[16]), .b(L15[10]), .cin(C15[9]), .f(L16[9]), .cout(C16[9]));
    adder_1 adder16_10(.a(X[10] & Y[16]), .b(L15[11]), .cin(C15[10]), .f(L16[10]), .cout(C16[10]));
    adder_1 adder16_11(.a(X[11] & Y[16]), .b(L15[12]), .cin(C15[11]), .f(L16[11]), .cout(C16[11]));
    adder_1 adder16_12(.a(X[12] & Y[16]), .b(L15[13]), .cin(C15[12]), .f(L16[12]), .cout(C16[12]));
    adder_1 adder16_13(.a(X[13] & Y[16]), .b(L15[14]), .cin(C15[13]), .f(L16[13]), .cout(C16[13]));
    adder_1 adder16_14(.a(X[14] & Y[16]), .b(L15[15]), .cin(C15[14]), .f(L16[14]), .cout(C16[14]));
    adder_1 adder16_15(.a(X[15] & Y[16]), .b(L15[16]), .cin(C15[15]), .f(L16[15]), .cout(C16[15]));
    adder_1 adder16_16(.a(X[16] & Y[16]), .b(L15[17]), .cin(C15[16]), .f(L16[16]), .cout(C16[16]));
    adder_1 adder16_17(.a(X[17] & Y[16]), .b(L15[18]), .cin(C15[17]), .f(L16[17]), .cout(C16[17]));
    adder_1 adder16_18(.a(X[18] & Y[16]), .b(L15[19]), .cin(C15[18]), .f(L16[18]), .cout(C16[18]));
    adder_1 adder16_19(.a(X[19] & Y[16]), .b(L15[20]), .cin(C15[19]), .f(L16[19]), .cout(C16[19]));
    adder_1 adder16_20(.a(X[20] & Y[16]), .b(L15[21]), .cin(C15[20]), .f(L16[20]), .cout(C16[20]));
    adder_1 adder16_21(.a(X[21] & Y[16]), .b(L15[22]), .cin(C15[21]), .f(L16[21]), .cout(C16[21]));
    adder_1 adder16_22(.a(X[22] & Y[16]), .b(L15[23]), .cin(C15[22]), .f(L16[22]), .cout(C16[22]));
    adder_1 adder16_23(.a(X[23] & Y[16]), .b(L15[24]), .cin(C15[23]), .f(L16[23]), .cout(C16[23]));
    adder_1 adder16_24(.a(X[24] & Y[16]), .b(L15[25]), .cin(C15[24]), .f(L16[24]), .cout(C16[24]));
    adder_1 adder16_25(.a(X[25] & Y[16]), .b(L15[26]), .cin(C15[25]), .f(L16[25]), .cout(C16[25]));
    adder_1 adder16_26(.a(X[26] & Y[16]), .b(L15[27]), .cin(C15[26]), .f(L16[26]), .cout(C16[26]));
    adder_1 adder16_27(.a(X[27] & Y[16]), .b(L15[28]), .cin(C15[27]), .f(L16[27]), .cout(C16[27]));
    adder_1 adder16_28(.a(X[28] & Y[16]), .b(L15[29]), .cin(C15[28]), .f(L16[28]), .cout(C16[28]));
    adder_1 adder16_29(.a(X[29] & Y[16]), .b(L15[30]), .cin(C15[29]), .f(L16[29]), .cout(C16[29]));
    adder_1 adder16_30(.a(X[30] & Y[16]), .b(L15[31]), .cin(C15[30]), .f(L16[30]), .cout(C16[30]));
    assign L16[31] = X[31] & Y[16];
    wire [31:0] L17, C17;
    adder_1 adder17_0(.a(X[0] & Y[17]), .b(L16[1]), .cin(C16[0]), .f(L17[0]), .cout(C17[0]));
    adder_1 adder17_1(.a(X[1] & Y[17]), .b(L16[2]), .cin(C16[1]), .f(L17[1]), .cout(C17[1]));
    adder_1 adder17_2(.a(X[2] & Y[17]), .b(L16[3]), .cin(C16[2]), .f(L17[2]), .cout(C17[2]));
    adder_1 adder17_3(.a(X[3] & Y[17]), .b(L16[4]), .cin(C16[3]), .f(L17[3]), .cout(C17[3]));
    adder_1 adder17_4(.a(X[4] & Y[17]), .b(L16[5]), .cin(C16[4]), .f(L17[4]), .cout(C17[4]));
    adder_1 adder17_5(.a(X[5] & Y[17]), .b(L16[6]), .cin(C16[5]), .f(L17[5]), .cout(C17[5]));
    adder_1 adder17_6(.a(X[6] & Y[17]), .b(L16[7]), .cin(C16[6]), .f(L17[6]), .cout(C17[6]));
    adder_1 adder17_7(.a(X[7] & Y[17]), .b(L16[8]), .cin(C16[7]), .f(L17[7]), .cout(C17[7]));
    adder_1 adder17_8(.a(X[8] & Y[17]), .b(L16[9]), .cin(C16[8]), .f(L17[8]), .cout(C17[8]));
    adder_1 adder17_9(.a(X[9] & Y[17]), .b(L16[10]), .cin(C16[9]), .f(L17[9]), .cout(C17[9]));
    adder_1 adder17_10(.a(X[10] & Y[17]), .b(L16[11]), .cin(C16[10]), .f(L17[10]), .cout(C17[10]));
    adder_1 adder17_11(.a(X[11] & Y[17]), .b(L16[12]), .cin(C16[11]), .f(L17[11]), .cout(C17[11]));
    adder_1 adder17_12(.a(X[12] & Y[17]), .b(L16[13]), .cin(C16[12]), .f(L17[12]), .cout(C17[12]));
    adder_1 adder17_13(.a(X[13] & Y[17]), .b(L16[14]), .cin(C16[13]), .f(L17[13]), .cout(C17[13]));
    adder_1 adder17_14(.a(X[14] & Y[17]), .b(L16[15]), .cin(C16[14]), .f(L17[14]), .cout(C17[14]));
    adder_1 adder17_15(.a(X[15] & Y[17]), .b(L16[16]), .cin(C16[15]), .f(L17[15]), .cout(C17[15]));
    adder_1 adder17_16(.a(X[16] & Y[17]), .b(L16[17]), .cin(C16[16]), .f(L17[16]), .cout(C17[16]));
    adder_1 adder17_17(.a(X[17] & Y[17]), .b(L16[18]), .cin(C16[17]), .f(L17[17]), .cout(C17[17]));
    adder_1 adder17_18(.a(X[18] & Y[17]), .b(L16[19]), .cin(C16[18]), .f(L17[18]), .cout(C17[18]));
    adder_1 adder17_19(.a(X[19] & Y[17]), .b(L16[20]), .cin(C16[19]), .f(L17[19]), .cout(C17[19]));
    adder_1 adder17_20(.a(X[20] & Y[17]), .b(L16[21]), .cin(C16[20]), .f(L17[20]), .cout(C17[20]));
    adder_1 adder17_21(.a(X[21] & Y[17]), .b(L16[22]), .cin(C16[21]), .f(L17[21]), .cout(C17[21]));
    adder_1 adder17_22(.a(X[22] & Y[17]), .b(L16[23]), .cin(C16[22]), .f(L17[22]), .cout(C17[22]));
    adder_1 adder17_23(.a(X[23] & Y[17]), .b(L16[24]), .cin(C16[23]), .f(L17[23]), .cout(C17[23]));
    adder_1 adder17_24(.a(X[24] & Y[17]), .b(L16[25]), .cin(C16[24]), .f(L17[24]), .cout(C17[24]));
    adder_1 adder17_25(.a(X[25] & Y[17]), .b(L16[26]), .cin(C16[25]), .f(L17[25]), .cout(C17[25]));
    adder_1 adder17_26(.a(X[26] & Y[17]), .b(L16[27]), .cin(C16[26]), .f(L17[26]), .cout(C17[26]));
    adder_1 adder17_27(.a(X[27] & Y[17]), .b(L16[28]), .cin(C16[27]), .f(L17[27]), .cout(C17[27]));
    adder_1 adder17_28(.a(X[28] & Y[17]), .b(L16[29]), .cin(C16[28]), .f(L17[28]), .cout(C17[28]));
    adder_1 adder17_29(.a(X[29] & Y[17]), .b(L16[30]), .cin(C16[29]), .f(L17[29]), .cout(C17[29]));
    adder_1 adder17_30(.a(X[30] & Y[17]), .b(L16[31]), .cin(C16[30]), .f(L17[30]), .cout(C17[30]));
    assign L17[31] = X[31] & Y[17];
    wire [31:0] L18, C18;
    adder_1 adder18_0(.a(X[0] & Y[18]), .b(L17[1]), .cin(C17[0]), .f(L18[0]), .cout(C18[0]));
    adder_1 adder18_1(.a(X[1] & Y[18]), .b(L17[2]), .cin(C17[1]), .f(L18[1]), .cout(C18[1]));
    adder_1 adder18_2(.a(X[2] & Y[18]), .b(L17[3]), .cin(C17[2]), .f(L18[2]), .cout(C18[2]));
    adder_1 adder18_3(.a(X[3] & Y[18]), .b(L17[4]), .cin(C17[3]), .f(L18[3]), .cout(C18[3]));
    adder_1 adder18_4(.a(X[4] & Y[18]), .b(L17[5]), .cin(C17[4]), .f(L18[4]), .cout(C18[4]));
    adder_1 adder18_5(.a(X[5] & Y[18]), .b(L17[6]), .cin(C17[5]), .f(L18[5]), .cout(C18[5]));
    adder_1 adder18_6(.a(X[6] & Y[18]), .b(L17[7]), .cin(C17[6]), .f(L18[6]), .cout(C18[6]));
    adder_1 adder18_7(.a(X[7] & Y[18]), .b(L17[8]), .cin(C17[7]), .f(L18[7]), .cout(C18[7]));
    adder_1 adder18_8(.a(X[8] & Y[18]), .b(L17[9]), .cin(C17[8]), .f(L18[8]), .cout(C18[8]));
    adder_1 adder18_9(.a(X[9] & Y[18]), .b(L17[10]), .cin(C17[9]), .f(L18[9]), .cout(C18[9]));
    adder_1 adder18_10(.a(X[10] & Y[18]), .b(L17[11]), .cin(C17[10]), .f(L18[10]), .cout(C18[10]));
    adder_1 adder18_11(.a(X[11] & Y[18]), .b(L17[12]), .cin(C17[11]), .f(L18[11]), .cout(C18[11]));
    adder_1 adder18_12(.a(X[12] & Y[18]), .b(L17[13]), .cin(C17[12]), .f(L18[12]), .cout(C18[12]));
    adder_1 adder18_13(.a(X[13] & Y[18]), .b(L17[14]), .cin(C17[13]), .f(L18[13]), .cout(C18[13]));
    adder_1 adder18_14(.a(X[14] & Y[18]), .b(L17[15]), .cin(C17[14]), .f(L18[14]), .cout(C18[14]));
    adder_1 adder18_15(.a(X[15] & Y[18]), .b(L17[16]), .cin(C17[15]), .f(L18[15]), .cout(C18[15]));
    adder_1 adder18_16(.a(X[16] & Y[18]), .b(L17[17]), .cin(C17[16]), .f(L18[16]), .cout(C18[16]));
    adder_1 adder18_17(.a(X[17] & Y[18]), .b(L17[18]), .cin(C17[17]), .f(L18[17]), .cout(C18[17]));
    adder_1 adder18_18(.a(X[18] & Y[18]), .b(L17[19]), .cin(C17[18]), .f(L18[18]), .cout(C18[18]));
    adder_1 adder18_19(.a(X[19] & Y[18]), .b(L17[20]), .cin(C17[19]), .f(L18[19]), .cout(C18[19]));
    adder_1 adder18_20(.a(X[20] & Y[18]), .b(L17[21]), .cin(C17[20]), .f(L18[20]), .cout(C18[20]));
    adder_1 adder18_21(.a(X[21] & Y[18]), .b(L17[22]), .cin(C17[21]), .f(L18[21]), .cout(C18[21]));
    adder_1 adder18_22(.a(X[22] & Y[18]), .b(L17[23]), .cin(C17[22]), .f(L18[22]), .cout(C18[22]));
    adder_1 adder18_23(.a(X[23] & Y[18]), .b(L17[24]), .cin(C17[23]), .f(L18[23]), .cout(C18[23]));
    adder_1 adder18_24(.a(X[24] & Y[18]), .b(L17[25]), .cin(C17[24]), .f(L18[24]), .cout(C18[24]));
    adder_1 adder18_25(.a(X[25] & Y[18]), .b(L17[26]), .cin(C17[25]), .f(L18[25]), .cout(C18[25]));
    adder_1 adder18_26(.a(X[26] & Y[18]), .b(L17[27]), .cin(C17[26]), .f(L18[26]), .cout(C18[26]));
    adder_1 adder18_27(.a(X[27] & Y[18]), .b(L17[28]), .cin(C17[27]), .f(L18[27]), .cout(C18[27]));
    adder_1 adder18_28(.a(X[28] & Y[18]), .b(L17[29]), .cin(C17[28]), .f(L18[28]), .cout(C18[28]));
    adder_1 adder18_29(.a(X[29] & Y[18]), .b(L17[30]), .cin(C17[29]), .f(L18[29]), .cout(C18[29]));
    adder_1 adder18_30(.a(X[30] & Y[18]), .b(L17[31]), .cin(C17[30]), .f(L18[30]), .cout(C18[30]));
    assign L18[31] = X[31] & Y[18];
    wire [31:0] L19, C19;
    adder_1 adder19_0(.a(X[0] & Y[19]), .b(L18[1]), .cin(C18[0]), .f(L19[0]), .cout(C19[0]));
    adder_1 adder19_1(.a(X[1] & Y[19]), .b(L18[2]), .cin(C18[1]), .f(L19[1]), .cout(C19[1]));
    adder_1 adder19_2(.a(X[2] & Y[19]), .b(L18[3]), .cin(C18[2]), .f(L19[2]), .cout(C19[2]));
    adder_1 adder19_3(.a(X[3] & Y[19]), .b(L18[4]), .cin(C18[3]), .f(L19[3]), .cout(C19[3]));
    adder_1 adder19_4(.a(X[4] & Y[19]), .b(L18[5]), .cin(C18[4]), .f(L19[4]), .cout(C19[4]));
    adder_1 adder19_5(.a(X[5] & Y[19]), .b(L18[6]), .cin(C18[5]), .f(L19[5]), .cout(C19[5]));
    adder_1 adder19_6(.a(X[6] & Y[19]), .b(L18[7]), .cin(C18[6]), .f(L19[6]), .cout(C19[6]));
    adder_1 adder19_7(.a(X[7] & Y[19]), .b(L18[8]), .cin(C18[7]), .f(L19[7]), .cout(C19[7]));
    adder_1 adder19_8(.a(X[8] & Y[19]), .b(L18[9]), .cin(C18[8]), .f(L19[8]), .cout(C19[8]));
    adder_1 adder19_9(.a(X[9] & Y[19]), .b(L18[10]), .cin(C18[9]), .f(L19[9]), .cout(C19[9]));
    adder_1 adder19_10(.a(X[10] & Y[19]), .b(L18[11]), .cin(C18[10]), .f(L19[10]), .cout(C19[10]));
    adder_1 adder19_11(.a(X[11] & Y[19]), .b(L18[12]), .cin(C18[11]), .f(L19[11]), .cout(C19[11]));
    adder_1 adder19_12(.a(X[12] & Y[19]), .b(L18[13]), .cin(C18[12]), .f(L19[12]), .cout(C19[12]));
    adder_1 adder19_13(.a(X[13] & Y[19]), .b(L18[14]), .cin(C18[13]), .f(L19[13]), .cout(C19[13]));
    adder_1 adder19_14(.a(X[14] & Y[19]), .b(L18[15]), .cin(C18[14]), .f(L19[14]), .cout(C19[14]));
    adder_1 adder19_15(.a(X[15] & Y[19]), .b(L18[16]), .cin(C18[15]), .f(L19[15]), .cout(C19[15]));
    adder_1 adder19_16(.a(X[16] & Y[19]), .b(L18[17]), .cin(C18[16]), .f(L19[16]), .cout(C19[16]));
    adder_1 adder19_17(.a(X[17] & Y[19]), .b(L18[18]), .cin(C18[17]), .f(L19[17]), .cout(C19[17]));
    adder_1 adder19_18(.a(X[18] & Y[19]), .b(L18[19]), .cin(C18[18]), .f(L19[18]), .cout(C19[18]));
    adder_1 adder19_19(.a(X[19] & Y[19]), .b(L18[20]), .cin(C18[19]), .f(L19[19]), .cout(C19[19]));
    adder_1 adder19_20(.a(X[20] & Y[19]), .b(L18[21]), .cin(C18[20]), .f(L19[20]), .cout(C19[20]));
    adder_1 adder19_21(.a(X[21] & Y[19]), .b(L18[22]), .cin(C18[21]), .f(L19[21]), .cout(C19[21]));
    adder_1 adder19_22(.a(X[22] & Y[19]), .b(L18[23]), .cin(C18[22]), .f(L19[22]), .cout(C19[22]));
    adder_1 adder19_23(.a(X[23] & Y[19]), .b(L18[24]), .cin(C18[23]), .f(L19[23]), .cout(C19[23]));
    adder_1 adder19_24(.a(X[24] & Y[19]), .b(L18[25]), .cin(C18[24]), .f(L19[24]), .cout(C19[24]));
    adder_1 adder19_25(.a(X[25] & Y[19]), .b(L18[26]), .cin(C18[25]), .f(L19[25]), .cout(C19[25]));
    adder_1 adder19_26(.a(X[26] & Y[19]), .b(L18[27]), .cin(C18[26]), .f(L19[26]), .cout(C19[26]));
    adder_1 adder19_27(.a(X[27] & Y[19]), .b(L18[28]), .cin(C18[27]), .f(L19[27]), .cout(C19[27]));
    adder_1 adder19_28(.a(X[28] & Y[19]), .b(L18[29]), .cin(C18[28]), .f(L19[28]), .cout(C19[28]));
    adder_1 adder19_29(.a(X[29] & Y[19]), .b(L18[30]), .cin(C18[29]), .f(L19[29]), .cout(C19[29]));
    adder_1 adder19_30(.a(X[30] & Y[19]), .b(L18[31]), .cin(C18[30]), .f(L19[30]), .cout(C19[30]));
    assign L19[31] = X[31] & Y[19];
    wire [31:0] L20, C20;
    adder_1 adder20_0(.a(X[0] & Y[20]), .b(L19[1]), .cin(C19[0]), .f(L20[0]), .cout(C20[0]));
    adder_1 adder20_1(.a(X[1] & Y[20]), .b(L19[2]), .cin(C19[1]), .f(L20[1]), .cout(C20[1]));
    adder_1 adder20_2(.a(X[2] & Y[20]), .b(L19[3]), .cin(C19[2]), .f(L20[2]), .cout(C20[2]));
    adder_1 adder20_3(.a(X[3] & Y[20]), .b(L19[4]), .cin(C19[3]), .f(L20[3]), .cout(C20[3]));
    adder_1 adder20_4(.a(X[4] & Y[20]), .b(L19[5]), .cin(C19[4]), .f(L20[4]), .cout(C20[4]));
    adder_1 adder20_5(.a(X[5] & Y[20]), .b(L19[6]), .cin(C19[5]), .f(L20[5]), .cout(C20[5]));
    adder_1 adder20_6(.a(X[6] & Y[20]), .b(L19[7]), .cin(C19[6]), .f(L20[6]), .cout(C20[6]));
    adder_1 adder20_7(.a(X[7] & Y[20]), .b(L19[8]), .cin(C19[7]), .f(L20[7]), .cout(C20[7]));
    adder_1 adder20_8(.a(X[8] & Y[20]), .b(L19[9]), .cin(C19[8]), .f(L20[8]), .cout(C20[8]));
    adder_1 adder20_9(.a(X[9] & Y[20]), .b(L19[10]), .cin(C19[9]), .f(L20[9]), .cout(C20[9]));
    adder_1 adder20_10(.a(X[10] & Y[20]), .b(L19[11]), .cin(C19[10]), .f(L20[10]), .cout(C20[10]));
    adder_1 adder20_11(.a(X[11] & Y[20]), .b(L19[12]), .cin(C19[11]), .f(L20[11]), .cout(C20[11]));
    adder_1 adder20_12(.a(X[12] & Y[20]), .b(L19[13]), .cin(C19[12]), .f(L20[12]), .cout(C20[12]));
    adder_1 adder20_13(.a(X[13] & Y[20]), .b(L19[14]), .cin(C19[13]), .f(L20[13]), .cout(C20[13]));
    adder_1 adder20_14(.a(X[14] & Y[20]), .b(L19[15]), .cin(C19[14]), .f(L20[14]), .cout(C20[14]));
    adder_1 adder20_15(.a(X[15] & Y[20]), .b(L19[16]), .cin(C19[15]), .f(L20[15]), .cout(C20[15]));
    adder_1 adder20_16(.a(X[16] & Y[20]), .b(L19[17]), .cin(C19[16]), .f(L20[16]), .cout(C20[16]));
    adder_1 adder20_17(.a(X[17] & Y[20]), .b(L19[18]), .cin(C19[17]), .f(L20[17]), .cout(C20[17]));
    adder_1 adder20_18(.a(X[18] & Y[20]), .b(L19[19]), .cin(C19[18]), .f(L20[18]), .cout(C20[18]));
    adder_1 adder20_19(.a(X[19] & Y[20]), .b(L19[20]), .cin(C19[19]), .f(L20[19]), .cout(C20[19]));
    adder_1 adder20_20(.a(X[20] & Y[20]), .b(L19[21]), .cin(C19[20]), .f(L20[20]), .cout(C20[20]));
    adder_1 adder20_21(.a(X[21] & Y[20]), .b(L19[22]), .cin(C19[21]), .f(L20[21]), .cout(C20[21]));
    adder_1 adder20_22(.a(X[22] & Y[20]), .b(L19[23]), .cin(C19[22]), .f(L20[22]), .cout(C20[22]));
    adder_1 adder20_23(.a(X[23] & Y[20]), .b(L19[24]), .cin(C19[23]), .f(L20[23]), .cout(C20[23]));
    adder_1 adder20_24(.a(X[24] & Y[20]), .b(L19[25]), .cin(C19[24]), .f(L20[24]), .cout(C20[24]));
    adder_1 adder20_25(.a(X[25] & Y[20]), .b(L19[26]), .cin(C19[25]), .f(L20[25]), .cout(C20[25]));
    adder_1 adder20_26(.a(X[26] & Y[20]), .b(L19[27]), .cin(C19[26]), .f(L20[26]), .cout(C20[26]));
    adder_1 adder20_27(.a(X[27] & Y[20]), .b(L19[28]), .cin(C19[27]), .f(L20[27]), .cout(C20[27]));
    adder_1 adder20_28(.a(X[28] & Y[20]), .b(L19[29]), .cin(C19[28]), .f(L20[28]), .cout(C20[28]));
    adder_1 adder20_29(.a(X[29] & Y[20]), .b(L19[30]), .cin(C19[29]), .f(L20[29]), .cout(C20[29]));
    adder_1 adder20_30(.a(X[30] & Y[20]), .b(L19[31]), .cin(C19[30]), .f(L20[30]), .cout(C20[30]));
    assign L20[31] = X[31] & Y[20];
    wire [31:0] L21, C21;
    adder_1 adder21_0(.a(X[0] & Y[21]), .b(L20[1]), .cin(C20[0]), .f(L21[0]), .cout(C21[0]));
    adder_1 adder21_1(.a(X[1] & Y[21]), .b(L20[2]), .cin(C20[1]), .f(L21[1]), .cout(C21[1]));
    adder_1 adder21_2(.a(X[2] & Y[21]), .b(L20[3]), .cin(C20[2]), .f(L21[2]), .cout(C21[2]));
    adder_1 adder21_3(.a(X[3] & Y[21]), .b(L20[4]), .cin(C20[3]), .f(L21[3]), .cout(C21[3]));
    adder_1 adder21_4(.a(X[4] & Y[21]), .b(L20[5]), .cin(C20[4]), .f(L21[4]), .cout(C21[4]));
    adder_1 adder21_5(.a(X[5] & Y[21]), .b(L20[6]), .cin(C20[5]), .f(L21[5]), .cout(C21[5]));
    adder_1 adder21_6(.a(X[6] & Y[21]), .b(L20[7]), .cin(C20[6]), .f(L21[6]), .cout(C21[6]));
    adder_1 adder21_7(.a(X[7] & Y[21]), .b(L20[8]), .cin(C20[7]), .f(L21[7]), .cout(C21[7]));
    adder_1 adder21_8(.a(X[8] & Y[21]), .b(L20[9]), .cin(C20[8]), .f(L21[8]), .cout(C21[8]));
    adder_1 adder21_9(.a(X[9] & Y[21]), .b(L20[10]), .cin(C20[9]), .f(L21[9]), .cout(C21[9]));
    adder_1 adder21_10(.a(X[10] & Y[21]), .b(L20[11]), .cin(C20[10]), .f(L21[10]), .cout(C21[10]));
    adder_1 adder21_11(.a(X[11] & Y[21]), .b(L20[12]), .cin(C20[11]), .f(L21[11]), .cout(C21[11]));
    adder_1 adder21_12(.a(X[12] & Y[21]), .b(L20[13]), .cin(C20[12]), .f(L21[12]), .cout(C21[12]));
    adder_1 adder21_13(.a(X[13] & Y[21]), .b(L20[14]), .cin(C20[13]), .f(L21[13]), .cout(C21[13]));
    adder_1 adder21_14(.a(X[14] & Y[21]), .b(L20[15]), .cin(C20[14]), .f(L21[14]), .cout(C21[14]));
    adder_1 adder21_15(.a(X[15] & Y[21]), .b(L20[16]), .cin(C20[15]), .f(L21[15]), .cout(C21[15]));
    adder_1 adder21_16(.a(X[16] & Y[21]), .b(L20[17]), .cin(C20[16]), .f(L21[16]), .cout(C21[16]));
    adder_1 adder21_17(.a(X[17] & Y[21]), .b(L20[18]), .cin(C20[17]), .f(L21[17]), .cout(C21[17]));
    adder_1 adder21_18(.a(X[18] & Y[21]), .b(L20[19]), .cin(C20[18]), .f(L21[18]), .cout(C21[18]));
    adder_1 adder21_19(.a(X[19] & Y[21]), .b(L20[20]), .cin(C20[19]), .f(L21[19]), .cout(C21[19]));
    adder_1 adder21_20(.a(X[20] & Y[21]), .b(L20[21]), .cin(C20[20]), .f(L21[20]), .cout(C21[20]));
    adder_1 adder21_21(.a(X[21] & Y[21]), .b(L20[22]), .cin(C20[21]), .f(L21[21]), .cout(C21[21]));
    adder_1 adder21_22(.a(X[22] & Y[21]), .b(L20[23]), .cin(C20[22]), .f(L21[22]), .cout(C21[22]));
    adder_1 adder21_23(.a(X[23] & Y[21]), .b(L20[24]), .cin(C20[23]), .f(L21[23]), .cout(C21[23]));
    adder_1 adder21_24(.a(X[24] & Y[21]), .b(L20[25]), .cin(C20[24]), .f(L21[24]), .cout(C21[24]));
    adder_1 adder21_25(.a(X[25] & Y[21]), .b(L20[26]), .cin(C20[25]), .f(L21[25]), .cout(C21[25]));
    adder_1 adder21_26(.a(X[26] & Y[21]), .b(L20[27]), .cin(C20[26]), .f(L21[26]), .cout(C21[26]));
    adder_1 adder21_27(.a(X[27] & Y[21]), .b(L20[28]), .cin(C20[27]), .f(L21[27]), .cout(C21[27]));
    adder_1 adder21_28(.a(X[28] & Y[21]), .b(L20[29]), .cin(C20[28]), .f(L21[28]), .cout(C21[28]));
    adder_1 adder21_29(.a(X[29] & Y[21]), .b(L20[30]), .cin(C20[29]), .f(L21[29]), .cout(C21[29]));
    adder_1 adder21_30(.a(X[30] & Y[21]), .b(L20[31]), .cin(C20[30]), .f(L21[30]), .cout(C21[30]));
    assign L21[31] = X[31] & Y[21];
    wire [31:0] L22, C22;
    adder_1 adder22_0(.a(X[0] & Y[22]), .b(L21[1]), .cin(C21[0]), .f(L22[0]), .cout(C22[0]));
    adder_1 adder22_1(.a(X[1] & Y[22]), .b(L21[2]), .cin(C21[1]), .f(L22[1]), .cout(C22[1]));
    adder_1 adder22_2(.a(X[2] & Y[22]), .b(L21[3]), .cin(C21[2]), .f(L22[2]), .cout(C22[2]));
    adder_1 adder22_3(.a(X[3] & Y[22]), .b(L21[4]), .cin(C21[3]), .f(L22[3]), .cout(C22[3]));
    adder_1 adder22_4(.a(X[4] & Y[22]), .b(L21[5]), .cin(C21[4]), .f(L22[4]), .cout(C22[4]));
    adder_1 adder22_5(.a(X[5] & Y[22]), .b(L21[6]), .cin(C21[5]), .f(L22[5]), .cout(C22[5]));
    adder_1 adder22_6(.a(X[6] & Y[22]), .b(L21[7]), .cin(C21[6]), .f(L22[6]), .cout(C22[6]));
    adder_1 adder22_7(.a(X[7] & Y[22]), .b(L21[8]), .cin(C21[7]), .f(L22[7]), .cout(C22[7]));
    adder_1 adder22_8(.a(X[8] & Y[22]), .b(L21[9]), .cin(C21[8]), .f(L22[8]), .cout(C22[8]));
    adder_1 adder22_9(.a(X[9] & Y[22]), .b(L21[10]), .cin(C21[9]), .f(L22[9]), .cout(C22[9]));
    adder_1 adder22_10(.a(X[10] & Y[22]), .b(L21[11]), .cin(C21[10]), .f(L22[10]), .cout(C22[10]));
    adder_1 adder22_11(.a(X[11] & Y[22]), .b(L21[12]), .cin(C21[11]), .f(L22[11]), .cout(C22[11]));
    adder_1 adder22_12(.a(X[12] & Y[22]), .b(L21[13]), .cin(C21[12]), .f(L22[12]), .cout(C22[12]));
    adder_1 adder22_13(.a(X[13] & Y[22]), .b(L21[14]), .cin(C21[13]), .f(L22[13]), .cout(C22[13]));
    adder_1 adder22_14(.a(X[14] & Y[22]), .b(L21[15]), .cin(C21[14]), .f(L22[14]), .cout(C22[14]));
    adder_1 adder22_15(.a(X[15] & Y[22]), .b(L21[16]), .cin(C21[15]), .f(L22[15]), .cout(C22[15]));
    adder_1 adder22_16(.a(X[16] & Y[22]), .b(L21[17]), .cin(C21[16]), .f(L22[16]), .cout(C22[16]));
    adder_1 adder22_17(.a(X[17] & Y[22]), .b(L21[18]), .cin(C21[17]), .f(L22[17]), .cout(C22[17]));
    adder_1 adder22_18(.a(X[18] & Y[22]), .b(L21[19]), .cin(C21[18]), .f(L22[18]), .cout(C22[18]));
    adder_1 adder22_19(.a(X[19] & Y[22]), .b(L21[20]), .cin(C21[19]), .f(L22[19]), .cout(C22[19]));
    adder_1 adder22_20(.a(X[20] & Y[22]), .b(L21[21]), .cin(C21[20]), .f(L22[20]), .cout(C22[20]));
    adder_1 adder22_21(.a(X[21] & Y[22]), .b(L21[22]), .cin(C21[21]), .f(L22[21]), .cout(C22[21]));
    adder_1 adder22_22(.a(X[22] & Y[22]), .b(L21[23]), .cin(C21[22]), .f(L22[22]), .cout(C22[22]));
    adder_1 adder22_23(.a(X[23] & Y[22]), .b(L21[24]), .cin(C21[23]), .f(L22[23]), .cout(C22[23]));
    adder_1 adder22_24(.a(X[24] & Y[22]), .b(L21[25]), .cin(C21[24]), .f(L22[24]), .cout(C22[24]));
    adder_1 adder22_25(.a(X[25] & Y[22]), .b(L21[26]), .cin(C21[25]), .f(L22[25]), .cout(C22[25]));
    adder_1 adder22_26(.a(X[26] & Y[22]), .b(L21[27]), .cin(C21[26]), .f(L22[26]), .cout(C22[26]));
    adder_1 adder22_27(.a(X[27] & Y[22]), .b(L21[28]), .cin(C21[27]), .f(L22[27]), .cout(C22[27]));
    adder_1 adder22_28(.a(X[28] & Y[22]), .b(L21[29]), .cin(C21[28]), .f(L22[28]), .cout(C22[28]));
    adder_1 adder22_29(.a(X[29] & Y[22]), .b(L21[30]), .cin(C21[29]), .f(L22[29]), .cout(C22[29]));
    adder_1 adder22_30(.a(X[30] & Y[22]), .b(L21[31]), .cin(C21[30]), .f(L22[30]), .cout(C22[30]));
    assign L22[31] = X[31] & Y[22];
    wire [31:0] L23, C23;
    adder_1 adder23_0(.a(X[0] & Y[23]), .b(L22[1]), .cin(C22[0]), .f(L23[0]), .cout(C23[0]));
    adder_1 adder23_1(.a(X[1] & Y[23]), .b(L22[2]), .cin(C22[1]), .f(L23[1]), .cout(C23[1]));
    adder_1 adder23_2(.a(X[2] & Y[23]), .b(L22[3]), .cin(C22[2]), .f(L23[2]), .cout(C23[2]));
    adder_1 adder23_3(.a(X[3] & Y[23]), .b(L22[4]), .cin(C22[3]), .f(L23[3]), .cout(C23[3]));
    adder_1 adder23_4(.a(X[4] & Y[23]), .b(L22[5]), .cin(C22[4]), .f(L23[4]), .cout(C23[4]));
    adder_1 adder23_5(.a(X[5] & Y[23]), .b(L22[6]), .cin(C22[5]), .f(L23[5]), .cout(C23[5]));
    adder_1 adder23_6(.a(X[6] & Y[23]), .b(L22[7]), .cin(C22[6]), .f(L23[6]), .cout(C23[6]));
    adder_1 adder23_7(.a(X[7] & Y[23]), .b(L22[8]), .cin(C22[7]), .f(L23[7]), .cout(C23[7]));
    adder_1 adder23_8(.a(X[8] & Y[23]), .b(L22[9]), .cin(C22[8]), .f(L23[8]), .cout(C23[8]));
    adder_1 adder23_9(.a(X[9] & Y[23]), .b(L22[10]), .cin(C22[9]), .f(L23[9]), .cout(C23[9]));
    adder_1 adder23_10(.a(X[10] & Y[23]), .b(L22[11]), .cin(C22[10]), .f(L23[10]), .cout(C23[10]));
    adder_1 adder23_11(.a(X[11] & Y[23]), .b(L22[12]), .cin(C22[11]), .f(L23[11]), .cout(C23[11]));
    adder_1 adder23_12(.a(X[12] & Y[23]), .b(L22[13]), .cin(C22[12]), .f(L23[12]), .cout(C23[12]));
    adder_1 adder23_13(.a(X[13] & Y[23]), .b(L22[14]), .cin(C22[13]), .f(L23[13]), .cout(C23[13]));
    adder_1 adder23_14(.a(X[14] & Y[23]), .b(L22[15]), .cin(C22[14]), .f(L23[14]), .cout(C23[14]));
    adder_1 adder23_15(.a(X[15] & Y[23]), .b(L22[16]), .cin(C22[15]), .f(L23[15]), .cout(C23[15]));
    adder_1 adder23_16(.a(X[16] & Y[23]), .b(L22[17]), .cin(C22[16]), .f(L23[16]), .cout(C23[16]));
    adder_1 adder23_17(.a(X[17] & Y[23]), .b(L22[18]), .cin(C22[17]), .f(L23[17]), .cout(C23[17]));
    adder_1 adder23_18(.a(X[18] & Y[23]), .b(L22[19]), .cin(C22[18]), .f(L23[18]), .cout(C23[18]));
    adder_1 adder23_19(.a(X[19] & Y[23]), .b(L22[20]), .cin(C22[19]), .f(L23[19]), .cout(C23[19]));
    adder_1 adder23_20(.a(X[20] & Y[23]), .b(L22[21]), .cin(C22[20]), .f(L23[20]), .cout(C23[20]));
    adder_1 adder23_21(.a(X[21] & Y[23]), .b(L22[22]), .cin(C22[21]), .f(L23[21]), .cout(C23[21]));
    adder_1 adder23_22(.a(X[22] & Y[23]), .b(L22[23]), .cin(C22[22]), .f(L23[22]), .cout(C23[22]));
    adder_1 adder23_23(.a(X[23] & Y[23]), .b(L22[24]), .cin(C22[23]), .f(L23[23]), .cout(C23[23]));
    adder_1 adder23_24(.a(X[24] & Y[23]), .b(L22[25]), .cin(C22[24]), .f(L23[24]), .cout(C23[24]));
    adder_1 adder23_25(.a(X[25] & Y[23]), .b(L22[26]), .cin(C22[25]), .f(L23[25]), .cout(C23[25]));
    adder_1 adder23_26(.a(X[26] & Y[23]), .b(L22[27]), .cin(C22[26]), .f(L23[26]), .cout(C23[26]));
    adder_1 adder23_27(.a(X[27] & Y[23]), .b(L22[28]), .cin(C22[27]), .f(L23[27]), .cout(C23[27]));
    adder_1 adder23_28(.a(X[28] & Y[23]), .b(L22[29]), .cin(C22[28]), .f(L23[28]), .cout(C23[28]));
    adder_1 adder23_29(.a(X[29] & Y[23]), .b(L22[30]), .cin(C22[29]), .f(L23[29]), .cout(C23[29]));
    adder_1 adder23_30(.a(X[30] & Y[23]), .b(L22[31]), .cin(C22[30]), .f(L23[30]), .cout(C23[30]));
    assign L23[31] = X[31] & Y[23];
    wire [31:0] L24, C24;
    adder_1 adder24_0(.a(X[0] & Y[24]), .b(L23[1]), .cin(C23[0]), .f(L24[0]), .cout(C24[0]));
    adder_1 adder24_1(.a(X[1] & Y[24]), .b(L23[2]), .cin(C23[1]), .f(L24[1]), .cout(C24[1]));
    adder_1 adder24_2(.a(X[2] & Y[24]), .b(L23[3]), .cin(C23[2]), .f(L24[2]), .cout(C24[2]));
    adder_1 adder24_3(.a(X[3] & Y[24]), .b(L23[4]), .cin(C23[3]), .f(L24[3]), .cout(C24[3]));
    adder_1 adder24_4(.a(X[4] & Y[24]), .b(L23[5]), .cin(C23[4]), .f(L24[4]), .cout(C24[4]));
    adder_1 adder24_5(.a(X[5] & Y[24]), .b(L23[6]), .cin(C23[5]), .f(L24[5]), .cout(C24[5]));
    adder_1 adder24_6(.a(X[6] & Y[24]), .b(L23[7]), .cin(C23[6]), .f(L24[6]), .cout(C24[6]));
    adder_1 adder24_7(.a(X[7] & Y[24]), .b(L23[8]), .cin(C23[7]), .f(L24[7]), .cout(C24[7]));
    adder_1 adder24_8(.a(X[8] & Y[24]), .b(L23[9]), .cin(C23[8]), .f(L24[8]), .cout(C24[8]));
    adder_1 adder24_9(.a(X[9] & Y[24]), .b(L23[10]), .cin(C23[9]), .f(L24[9]), .cout(C24[9]));
    adder_1 adder24_10(.a(X[10] & Y[24]), .b(L23[11]), .cin(C23[10]), .f(L24[10]), .cout(C24[10]));
    adder_1 adder24_11(.a(X[11] & Y[24]), .b(L23[12]), .cin(C23[11]), .f(L24[11]), .cout(C24[11]));
    adder_1 adder24_12(.a(X[12] & Y[24]), .b(L23[13]), .cin(C23[12]), .f(L24[12]), .cout(C24[12]));
    adder_1 adder24_13(.a(X[13] & Y[24]), .b(L23[14]), .cin(C23[13]), .f(L24[13]), .cout(C24[13]));
    adder_1 adder24_14(.a(X[14] & Y[24]), .b(L23[15]), .cin(C23[14]), .f(L24[14]), .cout(C24[14]));
    adder_1 adder24_15(.a(X[15] & Y[24]), .b(L23[16]), .cin(C23[15]), .f(L24[15]), .cout(C24[15]));
    adder_1 adder24_16(.a(X[16] & Y[24]), .b(L23[17]), .cin(C23[16]), .f(L24[16]), .cout(C24[16]));
    adder_1 adder24_17(.a(X[17] & Y[24]), .b(L23[18]), .cin(C23[17]), .f(L24[17]), .cout(C24[17]));
    adder_1 adder24_18(.a(X[18] & Y[24]), .b(L23[19]), .cin(C23[18]), .f(L24[18]), .cout(C24[18]));
    adder_1 adder24_19(.a(X[19] & Y[24]), .b(L23[20]), .cin(C23[19]), .f(L24[19]), .cout(C24[19]));
    adder_1 adder24_20(.a(X[20] & Y[24]), .b(L23[21]), .cin(C23[20]), .f(L24[20]), .cout(C24[20]));
    adder_1 adder24_21(.a(X[21] & Y[24]), .b(L23[22]), .cin(C23[21]), .f(L24[21]), .cout(C24[21]));
    adder_1 adder24_22(.a(X[22] & Y[24]), .b(L23[23]), .cin(C23[22]), .f(L24[22]), .cout(C24[22]));
    adder_1 adder24_23(.a(X[23] & Y[24]), .b(L23[24]), .cin(C23[23]), .f(L24[23]), .cout(C24[23]));
    adder_1 adder24_24(.a(X[24] & Y[24]), .b(L23[25]), .cin(C23[24]), .f(L24[24]), .cout(C24[24]));
    adder_1 adder24_25(.a(X[25] & Y[24]), .b(L23[26]), .cin(C23[25]), .f(L24[25]), .cout(C24[25]));
    adder_1 adder24_26(.a(X[26] & Y[24]), .b(L23[27]), .cin(C23[26]), .f(L24[26]), .cout(C24[26]));
    adder_1 adder24_27(.a(X[27] & Y[24]), .b(L23[28]), .cin(C23[27]), .f(L24[27]), .cout(C24[27]));
    adder_1 adder24_28(.a(X[28] & Y[24]), .b(L23[29]), .cin(C23[28]), .f(L24[28]), .cout(C24[28]));
    adder_1 adder24_29(.a(X[29] & Y[24]), .b(L23[30]), .cin(C23[29]), .f(L24[29]), .cout(C24[29]));
    adder_1 adder24_30(.a(X[30] & Y[24]), .b(L23[31]), .cin(C23[30]), .f(L24[30]), .cout(C24[30]));
    assign L24[31] = X[31] & Y[24];
    wire [31:0] L25, C25;
    adder_1 adder25_0(.a(X[0] & Y[25]), .b(L24[1]), .cin(C24[0]), .f(L25[0]), .cout(C25[0]));
    adder_1 adder25_1(.a(X[1] & Y[25]), .b(L24[2]), .cin(C24[1]), .f(L25[1]), .cout(C25[1]));
    adder_1 adder25_2(.a(X[2] & Y[25]), .b(L24[3]), .cin(C24[2]), .f(L25[2]), .cout(C25[2]));
    adder_1 adder25_3(.a(X[3] & Y[25]), .b(L24[4]), .cin(C24[3]), .f(L25[3]), .cout(C25[3]));
    adder_1 adder25_4(.a(X[4] & Y[25]), .b(L24[5]), .cin(C24[4]), .f(L25[4]), .cout(C25[4]));
    adder_1 adder25_5(.a(X[5] & Y[25]), .b(L24[6]), .cin(C24[5]), .f(L25[5]), .cout(C25[5]));
    adder_1 adder25_6(.a(X[6] & Y[25]), .b(L24[7]), .cin(C24[6]), .f(L25[6]), .cout(C25[6]));
    adder_1 adder25_7(.a(X[7] & Y[25]), .b(L24[8]), .cin(C24[7]), .f(L25[7]), .cout(C25[7]));
    adder_1 adder25_8(.a(X[8] & Y[25]), .b(L24[9]), .cin(C24[8]), .f(L25[8]), .cout(C25[8]));
    adder_1 adder25_9(.a(X[9] & Y[25]), .b(L24[10]), .cin(C24[9]), .f(L25[9]), .cout(C25[9]));
    adder_1 adder25_10(.a(X[10] & Y[25]), .b(L24[11]), .cin(C24[10]), .f(L25[10]), .cout(C25[10]));
    adder_1 adder25_11(.a(X[11] & Y[25]), .b(L24[12]), .cin(C24[11]), .f(L25[11]), .cout(C25[11]));
    adder_1 adder25_12(.a(X[12] & Y[25]), .b(L24[13]), .cin(C24[12]), .f(L25[12]), .cout(C25[12]));
    adder_1 adder25_13(.a(X[13] & Y[25]), .b(L24[14]), .cin(C24[13]), .f(L25[13]), .cout(C25[13]));
    adder_1 adder25_14(.a(X[14] & Y[25]), .b(L24[15]), .cin(C24[14]), .f(L25[14]), .cout(C25[14]));
    adder_1 adder25_15(.a(X[15] & Y[25]), .b(L24[16]), .cin(C24[15]), .f(L25[15]), .cout(C25[15]));
    adder_1 adder25_16(.a(X[16] & Y[25]), .b(L24[17]), .cin(C24[16]), .f(L25[16]), .cout(C25[16]));
    adder_1 adder25_17(.a(X[17] & Y[25]), .b(L24[18]), .cin(C24[17]), .f(L25[17]), .cout(C25[17]));
    adder_1 adder25_18(.a(X[18] & Y[25]), .b(L24[19]), .cin(C24[18]), .f(L25[18]), .cout(C25[18]));
    adder_1 adder25_19(.a(X[19] & Y[25]), .b(L24[20]), .cin(C24[19]), .f(L25[19]), .cout(C25[19]));
    adder_1 adder25_20(.a(X[20] & Y[25]), .b(L24[21]), .cin(C24[20]), .f(L25[20]), .cout(C25[20]));
    adder_1 adder25_21(.a(X[21] & Y[25]), .b(L24[22]), .cin(C24[21]), .f(L25[21]), .cout(C25[21]));
    adder_1 adder25_22(.a(X[22] & Y[25]), .b(L24[23]), .cin(C24[22]), .f(L25[22]), .cout(C25[22]));
    adder_1 adder25_23(.a(X[23] & Y[25]), .b(L24[24]), .cin(C24[23]), .f(L25[23]), .cout(C25[23]));
    adder_1 adder25_24(.a(X[24] & Y[25]), .b(L24[25]), .cin(C24[24]), .f(L25[24]), .cout(C25[24]));
    adder_1 adder25_25(.a(X[25] & Y[25]), .b(L24[26]), .cin(C24[25]), .f(L25[25]), .cout(C25[25]));
    adder_1 adder25_26(.a(X[26] & Y[25]), .b(L24[27]), .cin(C24[26]), .f(L25[26]), .cout(C25[26]));
    adder_1 adder25_27(.a(X[27] & Y[25]), .b(L24[28]), .cin(C24[27]), .f(L25[27]), .cout(C25[27]));
    adder_1 adder25_28(.a(X[28] & Y[25]), .b(L24[29]), .cin(C24[28]), .f(L25[28]), .cout(C25[28]));
    adder_1 adder25_29(.a(X[29] & Y[25]), .b(L24[30]), .cin(C24[29]), .f(L25[29]), .cout(C25[29]));
    adder_1 adder25_30(.a(X[30] & Y[25]), .b(L24[31]), .cin(C24[30]), .f(L25[30]), .cout(C25[30]));
    assign L25[31] = X[31] & Y[25];
    wire [31:0] L26, C26;
    adder_1 adder26_0(.a(X[0] & Y[26]), .b(L25[1]), .cin(C25[0]), .f(L26[0]), .cout(C26[0]));
    adder_1 adder26_1(.a(X[1] & Y[26]), .b(L25[2]), .cin(C25[1]), .f(L26[1]), .cout(C26[1]));
    adder_1 adder26_2(.a(X[2] & Y[26]), .b(L25[3]), .cin(C25[2]), .f(L26[2]), .cout(C26[2]));
    adder_1 adder26_3(.a(X[3] & Y[26]), .b(L25[4]), .cin(C25[3]), .f(L26[3]), .cout(C26[3]));
    adder_1 adder26_4(.a(X[4] & Y[26]), .b(L25[5]), .cin(C25[4]), .f(L26[4]), .cout(C26[4]));
    adder_1 adder26_5(.a(X[5] & Y[26]), .b(L25[6]), .cin(C25[5]), .f(L26[5]), .cout(C26[5]));
    adder_1 adder26_6(.a(X[6] & Y[26]), .b(L25[7]), .cin(C25[6]), .f(L26[6]), .cout(C26[6]));
    adder_1 adder26_7(.a(X[7] & Y[26]), .b(L25[8]), .cin(C25[7]), .f(L26[7]), .cout(C26[7]));
    adder_1 adder26_8(.a(X[8] & Y[26]), .b(L25[9]), .cin(C25[8]), .f(L26[8]), .cout(C26[8]));
    adder_1 adder26_9(.a(X[9] & Y[26]), .b(L25[10]), .cin(C25[9]), .f(L26[9]), .cout(C26[9]));
    adder_1 adder26_10(.a(X[10] & Y[26]), .b(L25[11]), .cin(C25[10]), .f(L26[10]), .cout(C26[10]));
    adder_1 adder26_11(.a(X[11] & Y[26]), .b(L25[12]), .cin(C25[11]), .f(L26[11]), .cout(C26[11]));
    adder_1 adder26_12(.a(X[12] & Y[26]), .b(L25[13]), .cin(C25[12]), .f(L26[12]), .cout(C26[12]));
    adder_1 adder26_13(.a(X[13] & Y[26]), .b(L25[14]), .cin(C25[13]), .f(L26[13]), .cout(C26[13]));
    adder_1 adder26_14(.a(X[14] & Y[26]), .b(L25[15]), .cin(C25[14]), .f(L26[14]), .cout(C26[14]));
    adder_1 adder26_15(.a(X[15] & Y[26]), .b(L25[16]), .cin(C25[15]), .f(L26[15]), .cout(C26[15]));
    adder_1 adder26_16(.a(X[16] & Y[26]), .b(L25[17]), .cin(C25[16]), .f(L26[16]), .cout(C26[16]));
    adder_1 adder26_17(.a(X[17] & Y[26]), .b(L25[18]), .cin(C25[17]), .f(L26[17]), .cout(C26[17]));
    adder_1 adder26_18(.a(X[18] & Y[26]), .b(L25[19]), .cin(C25[18]), .f(L26[18]), .cout(C26[18]));
    adder_1 adder26_19(.a(X[19] & Y[26]), .b(L25[20]), .cin(C25[19]), .f(L26[19]), .cout(C26[19]));
    adder_1 adder26_20(.a(X[20] & Y[26]), .b(L25[21]), .cin(C25[20]), .f(L26[20]), .cout(C26[20]));
    adder_1 adder26_21(.a(X[21] & Y[26]), .b(L25[22]), .cin(C25[21]), .f(L26[21]), .cout(C26[21]));
    adder_1 adder26_22(.a(X[22] & Y[26]), .b(L25[23]), .cin(C25[22]), .f(L26[22]), .cout(C26[22]));
    adder_1 adder26_23(.a(X[23] & Y[26]), .b(L25[24]), .cin(C25[23]), .f(L26[23]), .cout(C26[23]));
    adder_1 adder26_24(.a(X[24] & Y[26]), .b(L25[25]), .cin(C25[24]), .f(L26[24]), .cout(C26[24]));
    adder_1 adder26_25(.a(X[25] & Y[26]), .b(L25[26]), .cin(C25[25]), .f(L26[25]), .cout(C26[25]));
    adder_1 adder26_26(.a(X[26] & Y[26]), .b(L25[27]), .cin(C25[26]), .f(L26[26]), .cout(C26[26]));
    adder_1 adder26_27(.a(X[27] & Y[26]), .b(L25[28]), .cin(C25[27]), .f(L26[27]), .cout(C26[27]));
    adder_1 adder26_28(.a(X[28] & Y[26]), .b(L25[29]), .cin(C25[28]), .f(L26[28]), .cout(C26[28]));
    adder_1 adder26_29(.a(X[29] & Y[26]), .b(L25[30]), .cin(C25[29]), .f(L26[29]), .cout(C26[29]));
    adder_1 adder26_30(.a(X[30] & Y[26]), .b(L25[31]), .cin(C25[30]), .f(L26[30]), .cout(C26[30]));
    assign L26[31] = X[31] & Y[26];
    wire [31:0] L27, C27;
    adder_1 adder27_0(.a(X[0] & Y[27]), .b(L26[1]), .cin(C26[0]), .f(L27[0]), .cout(C27[0]));
    adder_1 adder27_1(.a(X[1] & Y[27]), .b(L26[2]), .cin(C26[1]), .f(L27[1]), .cout(C27[1]));
    adder_1 adder27_2(.a(X[2] & Y[27]), .b(L26[3]), .cin(C26[2]), .f(L27[2]), .cout(C27[2]));
    adder_1 adder27_3(.a(X[3] & Y[27]), .b(L26[4]), .cin(C26[3]), .f(L27[3]), .cout(C27[3]));
    adder_1 adder27_4(.a(X[4] & Y[27]), .b(L26[5]), .cin(C26[4]), .f(L27[4]), .cout(C27[4]));
    adder_1 adder27_5(.a(X[5] & Y[27]), .b(L26[6]), .cin(C26[5]), .f(L27[5]), .cout(C27[5]));
    adder_1 adder27_6(.a(X[6] & Y[27]), .b(L26[7]), .cin(C26[6]), .f(L27[6]), .cout(C27[6]));
    adder_1 adder27_7(.a(X[7] & Y[27]), .b(L26[8]), .cin(C26[7]), .f(L27[7]), .cout(C27[7]));
    adder_1 adder27_8(.a(X[8] & Y[27]), .b(L26[9]), .cin(C26[8]), .f(L27[8]), .cout(C27[8]));
    adder_1 adder27_9(.a(X[9] & Y[27]), .b(L26[10]), .cin(C26[9]), .f(L27[9]), .cout(C27[9]));
    adder_1 adder27_10(.a(X[10] & Y[27]), .b(L26[11]), .cin(C26[10]), .f(L27[10]), .cout(C27[10]));
    adder_1 adder27_11(.a(X[11] & Y[27]), .b(L26[12]), .cin(C26[11]), .f(L27[11]), .cout(C27[11]));
    adder_1 adder27_12(.a(X[12] & Y[27]), .b(L26[13]), .cin(C26[12]), .f(L27[12]), .cout(C27[12]));
    adder_1 adder27_13(.a(X[13] & Y[27]), .b(L26[14]), .cin(C26[13]), .f(L27[13]), .cout(C27[13]));
    adder_1 adder27_14(.a(X[14] & Y[27]), .b(L26[15]), .cin(C26[14]), .f(L27[14]), .cout(C27[14]));
    adder_1 adder27_15(.a(X[15] & Y[27]), .b(L26[16]), .cin(C26[15]), .f(L27[15]), .cout(C27[15]));
    adder_1 adder27_16(.a(X[16] & Y[27]), .b(L26[17]), .cin(C26[16]), .f(L27[16]), .cout(C27[16]));
    adder_1 adder27_17(.a(X[17] & Y[27]), .b(L26[18]), .cin(C26[17]), .f(L27[17]), .cout(C27[17]));
    adder_1 adder27_18(.a(X[18] & Y[27]), .b(L26[19]), .cin(C26[18]), .f(L27[18]), .cout(C27[18]));
    adder_1 adder27_19(.a(X[19] & Y[27]), .b(L26[20]), .cin(C26[19]), .f(L27[19]), .cout(C27[19]));
    adder_1 adder27_20(.a(X[20] & Y[27]), .b(L26[21]), .cin(C26[20]), .f(L27[20]), .cout(C27[20]));
    adder_1 adder27_21(.a(X[21] & Y[27]), .b(L26[22]), .cin(C26[21]), .f(L27[21]), .cout(C27[21]));
    adder_1 adder27_22(.a(X[22] & Y[27]), .b(L26[23]), .cin(C26[22]), .f(L27[22]), .cout(C27[22]));
    adder_1 adder27_23(.a(X[23] & Y[27]), .b(L26[24]), .cin(C26[23]), .f(L27[23]), .cout(C27[23]));
    adder_1 adder27_24(.a(X[24] & Y[27]), .b(L26[25]), .cin(C26[24]), .f(L27[24]), .cout(C27[24]));
    adder_1 adder27_25(.a(X[25] & Y[27]), .b(L26[26]), .cin(C26[25]), .f(L27[25]), .cout(C27[25]));
    adder_1 adder27_26(.a(X[26] & Y[27]), .b(L26[27]), .cin(C26[26]), .f(L27[26]), .cout(C27[26]));
    adder_1 adder27_27(.a(X[27] & Y[27]), .b(L26[28]), .cin(C26[27]), .f(L27[27]), .cout(C27[27]));
    adder_1 adder27_28(.a(X[28] & Y[27]), .b(L26[29]), .cin(C26[28]), .f(L27[28]), .cout(C27[28]));
    adder_1 adder27_29(.a(X[29] & Y[27]), .b(L26[30]), .cin(C26[29]), .f(L27[29]), .cout(C27[29]));
    adder_1 adder27_30(.a(X[30] & Y[27]), .b(L26[31]), .cin(C26[30]), .f(L27[30]), .cout(C27[30]));
    assign L27[31] = X[31] & Y[27];
    wire [31:0] L28, C28;
    adder_1 adder28_0(.a(X[0] & Y[28]), .b(L27[1]), .cin(C27[0]), .f(L28[0]), .cout(C28[0]));
    adder_1 adder28_1(.a(X[1] & Y[28]), .b(L27[2]), .cin(C27[1]), .f(L28[1]), .cout(C28[1]));
    adder_1 adder28_2(.a(X[2] & Y[28]), .b(L27[3]), .cin(C27[2]), .f(L28[2]), .cout(C28[2]));
    adder_1 adder28_3(.a(X[3] & Y[28]), .b(L27[4]), .cin(C27[3]), .f(L28[3]), .cout(C28[3]));
    adder_1 adder28_4(.a(X[4] & Y[28]), .b(L27[5]), .cin(C27[4]), .f(L28[4]), .cout(C28[4]));
    adder_1 adder28_5(.a(X[5] & Y[28]), .b(L27[6]), .cin(C27[5]), .f(L28[5]), .cout(C28[5]));
    adder_1 adder28_6(.a(X[6] & Y[28]), .b(L27[7]), .cin(C27[6]), .f(L28[6]), .cout(C28[6]));
    adder_1 adder28_7(.a(X[7] & Y[28]), .b(L27[8]), .cin(C27[7]), .f(L28[7]), .cout(C28[7]));
    adder_1 adder28_8(.a(X[8] & Y[28]), .b(L27[9]), .cin(C27[8]), .f(L28[8]), .cout(C28[8]));
    adder_1 adder28_9(.a(X[9] & Y[28]), .b(L27[10]), .cin(C27[9]), .f(L28[9]), .cout(C28[9]));
    adder_1 adder28_10(.a(X[10] & Y[28]), .b(L27[11]), .cin(C27[10]), .f(L28[10]), .cout(C28[10]));
    adder_1 adder28_11(.a(X[11] & Y[28]), .b(L27[12]), .cin(C27[11]), .f(L28[11]), .cout(C28[11]));
    adder_1 adder28_12(.a(X[12] & Y[28]), .b(L27[13]), .cin(C27[12]), .f(L28[12]), .cout(C28[12]));
    adder_1 adder28_13(.a(X[13] & Y[28]), .b(L27[14]), .cin(C27[13]), .f(L28[13]), .cout(C28[13]));
    adder_1 adder28_14(.a(X[14] & Y[28]), .b(L27[15]), .cin(C27[14]), .f(L28[14]), .cout(C28[14]));
    adder_1 adder28_15(.a(X[15] & Y[28]), .b(L27[16]), .cin(C27[15]), .f(L28[15]), .cout(C28[15]));
    adder_1 adder28_16(.a(X[16] & Y[28]), .b(L27[17]), .cin(C27[16]), .f(L28[16]), .cout(C28[16]));
    adder_1 adder28_17(.a(X[17] & Y[28]), .b(L27[18]), .cin(C27[17]), .f(L28[17]), .cout(C28[17]));
    adder_1 adder28_18(.a(X[18] & Y[28]), .b(L27[19]), .cin(C27[18]), .f(L28[18]), .cout(C28[18]));
    adder_1 adder28_19(.a(X[19] & Y[28]), .b(L27[20]), .cin(C27[19]), .f(L28[19]), .cout(C28[19]));
    adder_1 adder28_20(.a(X[20] & Y[28]), .b(L27[21]), .cin(C27[20]), .f(L28[20]), .cout(C28[20]));
    adder_1 adder28_21(.a(X[21] & Y[28]), .b(L27[22]), .cin(C27[21]), .f(L28[21]), .cout(C28[21]));
    adder_1 adder28_22(.a(X[22] & Y[28]), .b(L27[23]), .cin(C27[22]), .f(L28[22]), .cout(C28[22]));
    adder_1 adder28_23(.a(X[23] & Y[28]), .b(L27[24]), .cin(C27[23]), .f(L28[23]), .cout(C28[23]));
    adder_1 adder28_24(.a(X[24] & Y[28]), .b(L27[25]), .cin(C27[24]), .f(L28[24]), .cout(C28[24]));
    adder_1 adder28_25(.a(X[25] & Y[28]), .b(L27[26]), .cin(C27[25]), .f(L28[25]), .cout(C28[25]));
    adder_1 adder28_26(.a(X[26] & Y[28]), .b(L27[27]), .cin(C27[26]), .f(L28[26]), .cout(C28[26]));
    adder_1 adder28_27(.a(X[27] & Y[28]), .b(L27[28]), .cin(C27[27]), .f(L28[27]), .cout(C28[27]));
    adder_1 adder28_28(.a(X[28] & Y[28]), .b(L27[29]), .cin(C27[28]), .f(L28[28]), .cout(C28[28]));
    adder_1 adder28_29(.a(X[29] & Y[28]), .b(L27[30]), .cin(C27[29]), .f(L28[29]), .cout(C28[29]));
    adder_1 adder28_30(.a(X[30] & Y[28]), .b(L27[31]), .cin(C27[30]), .f(L28[30]), .cout(C28[30]));
    assign L28[31] = X[31] & Y[28];
    wire [31:0] L29, C29;
    adder_1 adder29_0(.a(X[0] & Y[29]), .b(L28[1]), .cin(C28[0]), .f(L29[0]), .cout(C29[0]));
    adder_1 adder29_1(.a(X[1] & Y[29]), .b(L28[2]), .cin(C28[1]), .f(L29[1]), .cout(C29[1]));
    adder_1 adder29_2(.a(X[2] & Y[29]), .b(L28[3]), .cin(C28[2]), .f(L29[2]), .cout(C29[2]));
    adder_1 adder29_3(.a(X[3] & Y[29]), .b(L28[4]), .cin(C28[3]), .f(L29[3]), .cout(C29[3]));
    adder_1 adder29_4(.a(X[4] & Y[29]), .b(L28[5]), .cin(C28[4]), .f(L29[4]), .cout(C29[4]));
    adder_1 adder29_5(.a(X[5] & Y[29]), .b(L28[6]), .cin(C28[5]), .f(L29[5]), .cout(C29[5]));
    adder_1 adder29_6(.a(X[6] & Y[29]), .b(L28[7]), .cin(C28[6]), .f(L29[6]), .cout(C29[6]));
    adder_1 adder29_7(.a(X[7] & Y[29]), .b(L28[8]), .cin(C28[7]), .f(L29[7]), .cout(C29[7]));
    adder_1 adder29_8(.a(X[8] & Y[29]), .b(L28[9]), .cin(C28[8]), .f(L29[8]), .cout(C29[8]));
    adder_1 adder29_9(.a(X[9] & Y[29]), .b(L28[10]), .cin(C28[9]), .f(L29[9]), .cout(C29[9]));
    adder_1 adder29_10(.a(X[10] & Y[29]), .b(L28[11]), .cin(C28[10]), .f(L29[10]), .cout(C29[10]));
    adder_1 adder29_11(.a(X[11] & Y[29]), .b(L28[12]), .cin(C28[11]), .f(L29[11]), .cout(C29[11]));
    adder_1 adder29_12(.a(X[12] & Y[29]), .b(L28[13]), .cin(C28[12]), .f(L29[12]), .cout(C29[12]));
    adder_1 adder29_13(.a(X[13] & Y[29]), .b(L28[14]), .cin(C28[13]), .f(L29[13]), .cout(C29[13]));
    adder_1 adder29_14(.a(X[14] & Y[29]), .b(L28[15]), .cin(C28[14]), .f(L29[14]), .cout(C29[14]));
    adder_1 adder29_15(.a(X[15] & Y[29]), .b(L28[16]), .cin(C28[15]), .f(L29[15]), .cout(C29[15]));
    adder_1 adder29_16(.a(X[16] & Y[29]), .b(L28[17]), .cin(C28[16]), .f(L29[16]), .cout(C29[16]));
    adder_1 adder29_17(.a(X[17] & Y[29]), .b(L28[18]), .cin(C28[17]), .f(L29[17]), .cout(C29[17]));
    adder_1 adder29_18(.a(X[18] & Y[29]), .b(L28[19]), .cin(C28[18]), .f(L29[18]), .cout(C29[18]));
    adder_1 adder29_19(.a(X[19] & Y[29]), .b(L28[20]), .cin(C28[19]), .f(L29[19]), .cout(C29[19]));
    adder_1 adder29_20(.a(X[20] & Y[29]), .b(L28[21]), .cin(C28[20]), .f(L29[20]), .cout(C29[20]));
    adder_1 adder29_21(.a(X[21] & Y[29]), .b(L28[22]), .cin(C28[21]), .f(L29[21]), .cout(C29[21]));
    adder_1 adder29_22(.a(X[22] & Y[29]), .b(L28[23]), .cin(C28[22]), .f(L29[22]), .cout(C29[22]));
    adder_1 adder29_23(.a(X[23] & Y[29]), .b(L28[24]), .cin(C28[23]), .f(L29[23]), .cout(C29[23]));
    adder_1 adder29_24(.a(X[24] & Y[29]), .b(L28[25]), .cin(C28[24]), .f(L29[24]), .cout(C29[24]));
    adder_1 adder29_25(.a(X[25] & Y[29]), .b(L28[26]), .cin(C28[25]), .f(L29[25]), .cout(C29[25]));
    adder_1 adder29_26(.a(X[26] & Y[29]), .b(L28[27]), .cin(C28[26]), .f(L29[26]), .cout(C29[26]));
    adder_1 adder29_27(.a(X[27] & Y[29]), .b(L28[28]), .cin(C28[27]), .f(L29[27]), .cout(C29[27]));
    adder_1 adder29_28(.a(X[28] & Y[29]), .b(L28[29]), .cin(C28[28]), .f(L29[28]), .cout(C29[28]));
    adder_1 adder29_29(.a(X[29] & Y[29]), .b(L28[30]), .cin(C28[29]), .f(L29[29]), .cout(C29[29]));
    adder_1 adder29_30(.a(X[30] & Y[29]), .b(L28[31]), .cin(C28[30]), .f(L29[30]), .cout(C29[30]));
    assign L29[31] = X[31] & Y[29];
    wire [31:0] L30, C30;
    adder_1 adder30_0(.a(X[0] & Y[30]), .b(L29[1]), .cin(C29[0]), .f(L30[0]), .cout(C30[0]));
    adder_1 adder30_1(.a(X[1] & Y[30]), .b(L29[2]), .cin(C29[1]), .f(L30[1]), .cout(C30[1]));
    adder_1 adder30_2(.a(X[2] & Y[30]), .b(L29[3]), .cin(C29[2]), .f(L30[2]), .cout(C30[2]));
    adder_1 adder30_3(.a(X[3] & Y[30]), .b(L29[4]), .cin(C29[3]), .f(L30[3]), .cout(C30[3]));
    adder_1 adder30_4(.a(X[4] & Y[30]), .b(L29[5]), .cin(C29[4]), .f(L30[4]), .cout(C30[4]));
    adder_1 adder30_5(.a(X[5] & Y[30]), .b(L29[6]), .cin(C29[5]), .f(L30[5]), .cout(C30[5]));
    adder_1 adder30_6(.a(X[6] & Y[30]), .b(L29[7]), .cin(C29[6]), .f(L30[6]), .cout(C30[6]));
    adder_1 adder30_7(.a(X[7] & Y[30]), .b(L29[8]), .cin(C29[7]), .f(L30[7]), .cout(C30[7]));
    adder_1 adder30_8(.a(X[8] & Y[30]), .b(L29[9]), .cin(C29[8]), .f(L30[8]), .cout(C30[8]));
    adder_1 adder30_9(.a(X[9] & Y[30]), .b(L29[10]), .cin(C29[9]), .f(L30[9]), .cout(C30[9]));
    adder_1 adder30_10(.a(X[10] & Y[30]), .b(L29[11]), .cin(C29[10]), .f(L30[10]), .cout(C30[10]));
    adder_1 adder30_11(.a(X[11] & Y[30]), .b(L29[12]), .cin(C29[11]), .f(L30[11]), .cout(C30[11]));
    adder_1 adder30_12(.a(X[12] & Y[30]), .b(L29[13]), .cin(C29[12]), .f(L30[12]), .cout(C30[12]));
    adder_1 adder30_13(.a(X[13] & Y[30]), .b(L29[14]), .cin(C29[13]), .f(L30[13]), .cout(C30[13]));
    adder_1 adder30_14(.a(X[14] & Y[30]), .b(L29[15]), .cin(C29[14]), .f(L30[14]), .cout(C30[14]));
    adder_1 adder30_15(.a(X[15] & Y[30]), .b(L29[16]), .cin(C29[15]), .f(L30[15]), .cout(C30[15]));
    adder_1 adder30_16(.a(X[16] & Y[30]), .b(L29[17]), .cin(C29[16]), .f(L30[16]), .cout(C30[16]));
    adder_1 adder30_17(.a(X[17] & Y[30]), .b(L29[18]), .cin(C29[17]), .f(L30[17]), .cout(C30[17]));
    adder_1 adder30_18(.a(X[18] & Y[30]), .b(L29[19]), .cin(C29[18]), .f(L30[18]), .cout(C30[18]));
    adder_1 adder30_19(.a(X[19] & Y[30]), .b(L29[20]), .cin(C29[19]), .f(L30[19]), .cout(C30[19]));
    adder_1 adder30_20(.a(X[20] & Y[30]), .b(L29[21]), .cin(C29[20]), .f(L30[20]), .cout(C30[20]));
    adder_1 adder30_21(.a(X[21] & Y[30]), .b(L29[22]), .cin(C29[21]), .f(L30[21]), .cout(C30[21]));
    adder_1 adder30_22(.a(X[22] & Y[30]), .b(L29[23]), .cin(C29[22]), .f(L30[22]), .cout(C30[22]));
    adder_1 adder30_23(.a(X[23] & Y[30]), .b(L29[24]), .cin(C29[23]), .f(L30[23]), .cout(C30[23]));
    adder_1 adder30_24(.a(X[24] & Y[30]), .b(L29[25]), .cin(C29[24]), .f(L30[24]), .cout(C30[24]));
    adder_1 adder30_25(.a(X[25] & Y[30]), .b(L29[26]), .cin(C29[25]), .f(L30[25]), .cout(C30[25]));
    adder_1 adder30_26(.a(X[26] & Y[30]), .b(L29[27]), .cin(C29[26]), .f(L30[26]), .cout(C30[26]));
    adder_1 adder30_27(.a(X[27] & Y[30]), .b(L29[28]), .cin(C29[27]), .f(L30[27]), .cout(C30[27]));
    adder_1 adder30_28(.a(X[28] & Y[30]), .b(L29[29]), .cin(C29[28]), .f(L30[28]), .cout(C30[28]));
    adder_1 adder30_29(.a(X[29] & Y[30]), .b(L29[30]), .cin(C29[29]), .f(L30[29]), .cout(C30[29]));
    adder_1 adder30_30(.a(X[30] & Y[30]), .b(L29[31]), .cin(C29[30]), .f(L30[30]), .cout(C30[30]));
    assign L30[31] = X[31] & Y[30];
    wire [31:0] L31, C31;
    adder_1 adder31_0(.a(X[0] & Y[31]), .b(L30[1]), .cin(C30[0]), .f(L31[0]), .cout(C31[0]));
    adder_1 adder31_1(.a(X[1] & Y[31]), .b(L30[2]), .cin(C30[1]), .f(L31[1]), .cout(C31[1]));
    adder_1 adder31_2(.a(X[2] & Y[31]), .b(L30[3]), .cin(C30[2]), .f(L31[2]), .cout(C31[2]));
    adder_1 adder31_3(.a(X[3] & Y[31]), .b(L30[4]), .cin(C30[3]), .f(L31[3]), .cout(C31[3]));
    adder_1 adder31_4(.a(X[4] & Y[31]), .b(L30[5]), .cin(C30[4]), .f(L31[4]), .cout(C31[4]));
    adder_1 adder31_5(.a(X[5] & Y[31]), .b(L30[6]), .cin(C30[5]), .f(L31[5]), .cout(C31[5]));
    adder_1 adder31_6(.a(X[6] & Y[31]), .b(L30[7]), .cin(C30[6]), .f(L31[6]), .cout(C31[6]));
    adder_1 adder31_7(.a(X[7] & Y[31]), .b(L30[8]), .cin(C30[7]), .f(L31[7]), .cout(C31[7]));
    adder_1 adder31_8(.a(X[8] & Y[31]), .b(L30[9]), .cin(C30[8]), .f(L31[8]), .cout(C31[8]));
    adder_1 adder31_9(.a(X[9] & Y[31]), .b(L30[10]), .cin(C30[9]), .f(L31[9]), .cout(C31[9]));
    adder_1 adder31_10(.a(X[10] & Y[31]), .b(L30[11]), .cin(C30[10]), .f(L31[10]), .cout(C31[10]));
    adder_1 adder31_11(.a(X[11] & Y[31]), .b(L30[12]), .cin(C30[11]), .f(L31[11]), .cout(C31[11]));
    adder_1 adder31_12(.a(X[12] & Y[31]), .b(L30[13]), .cin(C30[12]), .f(L31[12]), .cout(C31[12]));
    adder_1 adder31_13(.a(X[13] & Y[31]), .b(L30[14]), .cin(C30[13]), .f(L31[13]), .cout(C31[13]));
    adder_1 adder31_14(.a(X[14] & Y[31]), .b(L30[15]), .cin(C30[14]), .f(L31[14]), .cout(C31[14]));
    adder_1 adder31_15(.a(X[15] & Y[31]), .b(L30[16]), .cin(C30[15]), .f(L31[15]), .cout(C31[15]));
    adder_1 adder31_16(.a(X[16] & Y[31]), .b(L30[17]), .cin(C30[16]), .f(L31[16]), .cout(C31[16]));
    adder_1 adder31_17(.a(X[17] & Y[31]), .b(L30[18]), .cin(C30[17]), .f(L31[17]), .cout(C31[17]));
    adder_1 adder31_18(.a(X[18] & Y[31]), .b(L30[19]), .cin(C30[18]), .f(L31[18]), .cout(C31[18]));
    adder_1 adder31_19(.a(X[19] & Y[31]), .b(L30[20]), .cin(C30[19]), .f(L31[19]), .cout(C31[19]));
    adder_1 adder31_20(.a(X[20] & Y[31]), .b(L30[21]), .cin(C30[20]), .f(L31[20]), .cout(C31[20]));
    adder_1 adder31_21(.a(X[21] & Y[31]), .b(L30[22]), .cin(C30[21]), .f(L31[21]), .cout(C31[21]));
    adder_1 adder31_22(.a(X[22] & Y[31]), .b(L30[23]), .cin(C30[22]), .f(L31[22]), .cout(C31[22]));
    adder_1 adder31_23(.a(X[23] & Y[31]), .b(L30[24]), .cin(C30[23]), .f(L31[23]), .cout(C31[23]));
    adder_1 adder31_24(.a(X[24] & Y[31]), .b(L30[25]), .cin(C30[24]), .f(L31[24]), .cout(C31[24]));
    adder_1 adder31_25(.a(X[25] & Y[31]), .b(L30[26]), .cin(C30[25]), .f(L31[25]), .cout(C31[25]));
    adder_1 adder31_26(.a(X[26] & Y[31]), .b(L30[27]), .cin(C30[26]), .f(L31[26]), .cout(C31[26]));
    adder_1 adder31_27(.a(X[27] & Y[31]), .b(L30[28]), .cin(C30[27]), .f(L31[27]), .cout(C31[27]));
    adder_1 adder31_28(.a(X[28] & Y[31]), .b(L30[29]), .cin(C30[28]), .f(L31[28]), .cout(C31[28]));
    adder_1 adder31_29(.a(X[29] & Y[31]), .b(L30[30]), .cin(C30[29]), .f(L31[29]), .cout(C31[29]));
    adder_1 adder31_30(.a(X[30] & Y[31]), .b(L30[31]), .cin(C30[30]), .f(L31[30]), .cout(C31[30]));
    assign L31[31] = X[31] & Y[31];

    wire [31:0] L32, C32;
    /*
    ```python3
        for i in range(1, 31):
            print("adder_1 adder32_{}(.a(C31[{}]), .b(L31[{}]), .cin(C32[{}]), .f(L32[{}]), .cout(C32[{}]));".format(str(i), str(i), str(i+1), str(i-1), str(i), str(i)))
    ```
    */
    adder_1 adder32_0(.a(C31[0]), .b(L31[1]), .cin(1'b0), .f(L32[0]), .cout(C32[0]));
    adder_1 adder32_1(.a(C31[1]), .b(L31[2]), .cin(C32[0]), .f(L32[1]), .cout(C32[1]));
    adder_1 adder32_2(.a(C31[2]), .b(L31[3]), .cin(C32[1]), .f(L32[2]), .cout(C32[2]));
    adder_1 adder32_3(.a(C31[3]), .b(L31[4]), .cin(C32[2]), .f(L32[3]), .cout(C32[3]));
    adder_1 adder32_4(.a(C31[4]), .b(L31[5]), .cin(C32[3]), .f(L32[4]), .cout(C32[4]));
    adder_1 adder32_5(.a(C31[5]), .b(L31[6]), .cin(C32[4]), .f(L32[5]), .cout(C32[5]));
    adder_1 adder32_6(.a(C31[6]), .b(L31[7]), .cin(C32[5]), .f(L32[6]), .cout(C32[6]));
    adder_1 adder32_7(.a(C31[7]), .b(L31[8]), .cin(C32[6]), .f(L32[7]), .cout(C32[7]));
    adder_1 adder32_8(.a(C31[8]), .b(L31[9]), .cin(C32[7]), .f(L32[8]), .cout(C32[8]));
    adder_1 adder32_9(.a(C31[9]), .b(L31[10]), .cin(C32[8]), .f(L32[9]), .cout(C32[9]));
    adder_1 adder32_10(.a(C31[10]), .b(L31[11]), .cin(C32[9]), .f(L32[10]), .cout(C32[10]));
    adder_1 adder32_11(.a(C31[11]), .b(L31[12]), .cin(C32[10]), .f(L32[11]), .cout(C32[11]));
    adder_1 adder32_12(.a(C31[12]), .b(L31[13]), .cin(C32[11]), .f(L32[12]), .cout(C32[12]));
    adder_1 adder32_13(.a(C31[13]), .b(L31[14]), .cin(C32[12]), .f(L32[13]), .cout(C32[13]));
    adder_1 adder32_14(.a(C31[14]), .b(L31[15]), .cin(C32[13]), .f(L32[14]), .cout(C32[14]));
    adder_1 adder32_15(.a(C31[15]), .b(L31[16]), .cin(C32[14]), .f(L32[15]), .cout(C32[15]));
    adder_1 adder32_16(.a(C31[16]), .b(L31[17]), .cin(C32[15]), .f(L32[16]), .cout(C32[16]));
    adder_1 adder32_17(.a(C31[17]), .b(L31[18]), .cin(C32[16]), .f(L32[17]), .cout(C32[17]));
    adder_1 adder32_18(.a(C31[18]), .b(L31[19]), .cin(C32[17]), .f(L32[18]), .cout(C32[18]));
    adder_1 adder32_19(.a(C31[19]), .b(L31[20]), .cin(C32[18]), .f(L32[19]), .cout(C32[19]));
    adder_1 adder32_20(.a(C31[20]), .b(L31[21]), .cin(C32[19]), .f(L32[20]), .cout(C32[20]));
    adder_1 adder32_21(.a(C31[21]), .b(L31[22]), .cin(C32[20]), .f(L32[21]), .cout(C32[21]));
    adder_1 adder32_22(.a(C31[22]), .b(L31[23]), .cin(C32[21]), .f(L32[22]), .cout(C32[22]));
    adder_1 adder32_23(.a(C31[23]), .b(L31[24]), .cin(C32[22]), .f(L32[23]), .cout(C32[23]));
    adder_1 adder32_24(.a(C31[24]), .b(L31[25]), .cin(C32[23]), .f(L32[24]), .cout(C32[24]));
    adder_1 adder32_25(.a(C31[25]), .b(L31[26]), .cin(C32[24]), .f(L32[25]), .cout(C32[25]));
    adder_1 adder32_26(.a(C31[26]), .b(L31[27]), .cin(C32[25]), .f(L32[26]), .cout(C32[26]));
    adder_1 adder32_27(.a(C31[27]), .b(L31[28]), .cin(C32[26]), .f(L32[27]), .cout(C32[27]));
    adder_1 adder32_28(.a(C31[28]), .b(L31[29]), .cin(C32[27]), .f(L32[28]), .cout(C32[28]));
    adder_1 adder32_29(.a(C31[29]), .b(L31[30]), .cin(C32[28]), .f(L32[29]), .cout(C32[29]));
    adder_1 adder32_30(.a(C31[30]), .b(L31[31]), .cin(C32[29]), .f(L32[30]), .cout(C32[30]));
    assign L32[31] = C32[30];
    always @(*) begin
        /*
        ```python3
            for i in range(0, 32):
                print("P[{}] = L{}[0];".format(str(i), str(i)))
        ```
            */
        P[0] = L0[0];
        P[1] = L1[0];
        P[2] = L2[0];
        P[3] = L3[0];
        P[4] = L4[0];
        P[5] = L5[0];
        P[6] = L6[0];
        P[7] = L7[0];
        P[8] = L8[0];
        P[9] = L9[0];
        P[10] = L10[0];
        P[11] = L11[0];
        P[12] = L12[0];
        P[13] = L13[0];
        P[14] = L14[0];
        P[15] = L15[0];
        P[16] = L16[0];
        P[17] = L17[0];
        P[18] = L18[0];
        P[19] = L19[0];
        P[20] = L20[0];
        P[21] = L21[0];
        P[22] = L22[0];
        P[23] = L23[0];
        P[24] = L24[0];
        P[25] = L25[0];
        P[26] = L26[0];
        P[27] = L27[0];
        P[28] = L28[0];
        P[29] = L29[0];
        P[30] = L30[0];
        P[31] = L31[0];
        /*
        ```python3
            for i in range(0, 32):
                print("P[{}] = L32[{}];".format(str(32+i), str(i)))
        ```
        */
        P[32] = L32[0];
        P[33] = L32[1];
        P[34] = L32[2];
        P[35] = L32[3];
        P[36] = L32[4];
        P[37] = L32[5];
        P[38] = L32[6];
        P[39] = L32[7];
        P[40] = L32[8];
        P[41] = L32[9];
        P[42] = L32[10];
        P[43] = L32[11];
        P[44] = L32[12];
        P[45] = L32[13];
        P[46] = L32[14];
        P[47] = L32[15];
        P[48] = L32[16];
        P[49] = L32[17];
        P[50] = L32[18];
        P[51] = L32[19];
        P[52] = L32[20];
        P[53] = L32[21];
        P[54] = L32[22];
        P[55] = L32[23];
        P[56] = L32[24];
        P[57] = L32[25];
        P[58] = L32[26];
        P[59] = L32[27];
        P[60] = L32[28];
        P[61] = L32[29];
        P[62] = L32[30];
        P[63] = L32[31];
    end
endmodule
