
module term_man(
    input [31:0] addra,
    input [7:0] ascii_in,
    input [15:0] kbsig,//8:u, 7:d, 6:l, 5:r
    input clk,
    input in_valid,
    output [11:0] douta,
    output [2:0] state
);
    wire out;
    reg [7:0] text [2399:0];
    reg [31:0] ptr = 401;
    reg [2:0] state_R = 0;
    assign state = state_R;
    initial begin
        text[0] = 8'd45;
        text[1] = 8'd45;
        text[2] = 8'd45;
        text[3] = 8'd45;
        text[4] = 8'd45;
        text[5] = 8'd45;
        text[6] = 8'd45;
        text[7] = 8'd88;
        text[8] = 8'd116;
        text[9] = 8'd101;
        text[10] = 8'd114;
        text[11] = 8'd109;
        text[12] = 8'd105;
        text[13] = 8'd110;
        text[14] = 8'd97;
        text[15] = 8'd108;
        text[16] = 8'd45;
        text[17] = 8'd45;
        text[18] = 8'd45;
        text[19] = 8'd45;
        text[20] = 8'd45;
        text[21] = 8'd45;
        text[22] = 8'd45;
        text[23] = 8'd45;
        text[24] = 8'd45;
        text[25] = 8'd45;
        text[26] = 8'd45;
        text[27] = 8'd45;
        text[28] = 8'd45;
        text[29] = 8'd45;
        text[30] = 8'd45;
        text[31] = 8'd45;
        text[32] = 8'd45;
        text[33] = 8'd45;
        text[34] = 8'd45;
        text[35] = 8'd45;
        text[36] = 8'd45;
        text[37] = 8'd45;
        text[38] = 8'd45;
        text[39] = 8'd45;
        text[40] = 8'd45;
        text[41] = 8'd45;
        text[42] = 8'd91;
        text[43] = 8'd50;
        text[44] = 8'd49;
        text[45] = 8'd49;
        text[46] = 8'd53;
        text[47] = 8'd48;
        text[48] = 8'd50;
        text[49] = 8'd48;
        text[50] = 8'd48;
        text[51] = 8'd56;
        text[52] = 8'd93;
        text[53] = 8'd45;
        text[54] = 8'd45;
        text[55] = 8'd91;
        text[56] = 8'd67;
        text[57] = 8'd104;
        text[58] = 8'd101;
        text[59] = 8'd110;
        text[60] = 8'd103;
        text[61] = 8'd120;
        text[62] = 8'd105;
        text[63] = 8'd95;
        text[64] = 8'd76;
        text[65] = 8'd105;
        text[66] = 8'd93;
        text[67] = 8'd45;
        text[68] = 8'd45;
        text[69] = 8'd91;
        text[70] = 8'd50;
        text[71] = 8'd51;
        text[72] = 8'd58;
        text[73] = 8'd52;
        text[74] = 8'd58;
        text[75] = 8'd50;
        text[76] = 8'd51;
        text[77] = 8'd93;
        text[78] = 8'd45;
        text[79] = 8'd45;
        text[80] = 8'd91;
        text[81] = 8'd71;
        text[82] = 8'd93;
        text[83] = 8'd114;
        text[84] = 8'd97;
        text[85] = 8'd112;
        text[86] = 8'd104;
        text[87] = 8'd105;
        text[88] = 8'd99;
        text[89] = 8'd115;
        text[90] = 8'd32;
        text[91] = 8'd32;
        text[92] = 8'd32;
        text[93] = 8'd32;
        text[94] = 8'd32;
        text[95] = 8'd32;
        text[96] = 8'd32;
        text[97] = 8'd32;
        text[98] = 8'd32;
        text[99] = 8'd32;
        text[100] = 8'd32;
        text[101] = 8'd32;
        text[102] = 8'd32;
        text[103] = 8'd32;
        text[104] = 8'd32;
        text[105] = 8'd32;
        text[106] = 8'd32;
        text[107] = 8'd32;
        text[108] = 8'd32;
        text[109] = 8'd32;
        text[110] = 8'd32;
        text[111] = 8'd32;
        text[112] = 8'd32;
        text[113] = 8'd32;
        text[114] = 8'd32;
        text[115] = 8'd32;
        text[116] = 8'd32;
        text[117] = 8'd32;
        text[118] = 8'd32;
        text[119] = 8'd32;
        text[120] = 8'd32;
        text[121] = 8'd32;
        text[122] = 8'd32;
        text[123] = 8'd32;
        text[124] = 8'd32;
        text[125] = 8'd32;
        text[126] = 8'd32;
        text[127] = 8'd32;
        text[128] = 8'd32;
        text[129] = 8'd32;
        text[130] = 8'd32;
        text[131] = 8'd32;
        text[132] = 8'd32;
        text[133] = 8'd32;
        text[134] = 8'd32;
        text[135] = 8'd32;
        text[136] = 8'd32;
        text[137] = 8'd32;
        text[138] = 8'd32;
        text[139] = 8'd32;
        text[140] = 8'd32;
        text[141] = 8'd32;
        text[142] = 8'd32;
        text[143] = 8'd32;
        text[144] = 8'd32;
        text[145] = 8'd32;
        text[146] = 8'd32;
        text[147] = 8'd32;
        text[148] = 8'd32;
        text[149] = 8'd32;
        text[150] = 8'd32;
        text[151] = 8'd32;
        text[152] = 8'd32;
        text[153] = 8'd32;
        text[154] = 8'd32;
        text[155] = 8'd32;
        text[156] = 8'd32;
        text[157] = 8'd32;
        text[158] = 8'd32;
        text[159] = 8'd32;
        text[160] = 8'd91;
        text[161] = 8'd73;
        text[162] = 8'd93;
        text[163] = 8'd109;
        text[164] = 8'd97;
        text[165] = 8'd103;
        text[166] = 8'd101;
        text[167] = 8'd32;
        text[168] = 8'd32;
        text[169] = 8'd32;
        text[170] = 8'd32;
        text[171] = 8'd32;
        text[172] = 8'd32;
        text[173] = 8'd32;
        text[174] = 8'd32;
        text[175] = 8'd32;
        text[176] = 8'd32;
        text[177] = 8'd32;
        text[178] = 8'd32;
        text[179] = 8'd32;
        text[180] = 8'd32;
        text[181] = 8'd32;
        text[182] = 8'd32;
        text[183] = 8'd32;
        text[184] = 8'd32;
        text[185] = 8'd32;
        text[186] = 8'd32;
        text[187] = 8'd32;
        text[188] = 8'd32;
        text[189] = 8'd32;
        text[190] = 8'd32;
        text[191] = 8'd32;
        text[192] = 8'd32;
        text[193] = 8'd32;
        text[194] = 8'd32;
        text[195] = 8'd32;
        text[196] = 8'd32;
        text[197] = 8'd32;
        text[198] = 8'd32;
        text[199] = 8'd32;
        text[200] = 8'd32;
        text[201] = 8'd32;
        text[202] = 8'd32;
        text[203] = 8'd32;
        text[204] = 8'd32;
        text[205] = 8'd32;
        text[206] = 8'd32;
        text[207] = 8'd32;
        text[208] = 8'd32;
        text[209] = 8'd32;
        text[210] = 8'd32;
        text[211] = 8'd32;
        text[212] = 8'd32;
        text[213] = 8'd32;
        text[214] = 8'd32;
        text[215] = 8'd32;
        text[216] = 8'd32;
        text[217] = 8'd32;
        text[218] = 8'd32;
        text[219] = 8'd32;
        text[220] = 8'd32;
        text[221] = 8'd32;
        text[222] = 8'd32;
        text[223] = 8'd32;
        text[224] = 8'd32;
        text[225] = 8'd32;
        text[226] = 8'd32;
        text[227] = 8'd32;
        text[228] = 8'd32;
        text[229] = 8'd32;
        text[230] = 8'd32;
        text[231] = 8'd32;
        text[232] = 8'd32;
        text[233] = 8'd32;
        text[234] = 8'd32;
        text[235] = 8'd32;
        text[236] = 8'd32;
        text[237] = 8'd32;
        text[238] = 8'd32;
        text[239] = 8'd32;
        text[240] = 8'd91;
        text[241] = 8'd84;
        text[242] = 8'd93;
        text[243] = 8'd120;
        text[244] = 8'd116;
        text[245] = 8'd32;
        text[246] = 8'd32;
        text[247] = 8'd32;
        text[248] = 8'd32;
        text[249] = 8'd32;
        text[250] = 8'd32;
        text[251] = 8'd32;
        text[252] = 8'd32;
        text[253] = 8'd32;
        text[254] = 8'd32;
        text[255] = 8'd32;
        text[256] = 8'd32;
        text[257] = 8'd32;
        text[258] = 8'd32;
        text[259] = 8'd32;
        text[260] = 8'd32;
        text[261] = 8'd32;
        text[262] = 8'd32;
        text[263] = 8'd32;
        text[264] = 8'd32;
        text[265] = 8'd32;
        text[266] = 8'd32;
        text[267] = 8'd32;
        text[268] = 8'd32;
        text[269] = 8'd32;
        text[270] = 8'd32;
        text[271] = 8'd32;
        text[272] = 8'd32;
        text[273] = 8'd32;
        text[274] = 8'd32;
        text[275] = 8'd32;
        text[276] = 8'd32;
        text[277] = 8'd32;
        text[278] = 8'd32;
        text[279] = 8'd32;
        text[280] = 8'd32;
        text[281] = 8'd32;
        text[282] = 8'd32;
        text[283] = 8'd32;
        text[284] = 8'd32;
        text[285] = 8'd32;
        text[286] = 8'd32;
        text[287] = 8'd32;
        text[288] = 8'd32;
        text[289] = 8'd32;
        text[290] = 8'd32;
        text[291] = 8'd32;
        text[292] = 8'd32;
        text[293] = 8'd32;
        text[294] = 8'd32;
        text[295] = 8'd32;
        text[296] = 8'd32;
        text[297] = 8'd32;
        text[298] = 8'd32;
        text[299] = 8'd32;
        text[300] = 8'd32;
        text[301] = 8'd32;
        text[302] = 8'd32;
        text[303] = 8'd32;
        text[304] = 8'd32;
        text[305] = 8'd32;
        text[306] = 8'd32;
        text[307] = 8'd32;
        text[308] = 8'd32;
        text[309] = 8'd32;
        text[310] = 8'd32;
        text[311] = 8'd32;
        text[312] = 8'd32;
        text[313] = 8'd32;
        text[314] = 8'd32;
        text[315] = 8'd32;
        text[316] = 8'd32;
        text[317] = 8'd32;
        text[318] = 8'd32;
        text[319] = 8'd32;
        text[320] = 8'd91;
        text[321] = 8'd67;
        text[322] = 8'd93;
        text[323] = 8'd97;
        text[324] = 8'd108;
        text[325] = 8'd99;
        text[326] = 8'd117;
        text[327] = 8'd108;
        text[328] = 8'd97;
        text[329] = 8'd116;
        text[330] = 8'd111;
        text[331] = 8'd114;
        text[332] = 8'd32;
        text[333] = 8'd32;
        text[334] = 8'd32;
        text[335] = 8'd32;
        text[336] = 8'd32;
        text[337] = 8'd32;
        text[338] = 8'd32;
        text[339] = 8'd32;
        text[340] = 8'd32;
        text[341] = 8'd32;
        text[342] = 8'd32;
        text[343] = 8'd32;
        text[344] = 8'd32;
        text[345] = 8'd32;
        text[346] = 8'd32;
        text[347] = 8'd32;
        text[348] = 8'd32;
        text[349] = 8'd32;
        text[350] = 8'd32;
        text[351] = 8'd32;
        text[352] = 8'd32;
        text[353] = 8'd32;
        text[354] = 8'd32;
        text[355] = 8'd32;
        text[356] = 8'd32;
        text[357] = 8'd32;
        text[358] = 8'd32;
        text[359] = 8'd32;
        text[360] = 8'd32;
        text[361] = 8'd32;
        text[362] = 8'd32;
        text[363] = 8'd32;
        text[364] = 8'd32;
        text[365] = 8'd32;
        text[366] = 8'd32;
        text[367] = 8'd32;
        text[368] = 8'd32;
        text[369] = 8'd32;
        text[370] = 8'd32;
        text[371] = 8'd32;
        text[372] = 8'd32;
        text[373] = 8'd32;
        text[374] = 8'd32;
        text[375] = 8'd32;
        text[376] = 8'd32;
        text[377] = 8'd32;
        text[378] = 8'd32;
        text[379] = 8'd32;
        text[380] = 8'd32;
        text[381] = 8'd32;
        text[382] = 8'd32;
        text[383] = 8'd32;
        text[384] = 8'd32;
        text[385] = 8'd32;
        text[386] = 8'd32;
        text[387] = 8'd32;
        text[388] = 8'd32;
        text[389] = 8'd32;
        text[390] = 8'd32;
        text[391] = 8'd32;
        text[392] = 8'd32;
        text[393] = 8'd32;
        text[394] = 8'd32;
        text[395] = 8'd32;
        text[396] = 8'd32;
        text[397] = 8'd32;
        text[398] = 8'd32;
        text[399] = 8'd32;
        text[400] = 8'd45;
        text[401] = 8'd32;
        text[402] = 8'd32;
        text[403] = 8'd32;
        text[404] = 8'd32;
        text[405] = 8'd32;
        text[406] = 8'd32;
        text[407] = 8'd32;
        text[408] = 8'd32;
        text[409] = 8'd32;
        text[410] = 8'd32;
        text[411] = 8'd32;
        text[412] = 8'd32;
        text[413] = 8'd32;
        text[414] = 8'd32;
        text[415] = 8'd32;
        text[416] = 8'd32;
        text[417] = 8'd32;
        text[418] = 8'd32;
        text[419] = 8'd32;
        text[420] = 8'd32;
        text[421] = 8'd32;
        text[422] = 8'd32;
        text[423] = 8'd32;
        text[424] = 8'd32;
        text[425] = 8'd32;
        text[426] = 8'd32;
        text[427] = 8'd32;
        text[428] = 8'd32;
        text[429] = 8'd32;
        text[430] = 8'd32;
        text[431] = 8'd32;
        text[432] = 8'd32;
        text[433] = 8'd32;
        text[434] = 8'd32;
        text[435] = 8'd32;
        text[436] = 8'd32;
        text[437] = 8'd32;
        text[438] = 8'd32;
        text[439] = 8'd32;
        text[440] = 8'd32;
        text[441] = 8'd32;
        text[442] = 8'd32;
        text[443] = 8'd32;
        text[444] = 8'd32;
        text[445] = 8'd32;
        text[446] = 8'd32;
        text[447] = 8'd32;
        text[448] = 8'd32;
        text[449] = 8'd32;
        text[450] = 8'd32;
        text[451] = 8'd32;
        text[452] = 8'd32;
        text[453] = 8'd32;
        text[454] = 8'd32;
        text[455] = 8'd32;
        text[456] = 8'd32;
        text[457] = 8'd32;
        text[458] = 8'd32;
        text[459] = 8'd32;
        text[460] = 8'd32;
        text[461] = 8'd32;
        text[462] = 8'd32;
        text[463] = 8'd32;
        text[464] = 8'd32;
        text[465] = 8'd32;
        text[466] = 8'd32;
        text[467] = 8'd32;
        text[468] = 8'd32;
        text[469] = 8'd32;
        text[470] = 8'd32;
        text[471] = 8'd32;
        text[472] = 8'd32;
        text[473] = 8'd32;
        text[474] = 8'd32;
        text[475] = 8'd32;
        text[476] = 8'd32;
        text[477] = 8'd32;
        text[478] = 8'd32;
        text[479] = 8'd32;
    end
    wire [31:0] xw = addra % 8, yw = ((addra / 640) % 16);

    always @(posedge clk) begin
        if(kbsig[10] == 1) begin
            $display("ESC");
            state_R <= 0;
        end else if(state_R == 0) begin
            if(in_valid == 1) begin
                if(ascii_in == 8'h0D) begin
                    if(text[401] == 8'd84) begin
                        text[401] <= 0;
                        state_R <= 3;
                        ptr <= 32'd401;
                        $display("401 : %d", text[401]);
                        $display("state: %d", state_R);
                        text[480] = 8'd0;
                        text[481] = 8'd0;
                        text[482] = 8'd0;
                        text[483] = 8'd0;
                        text[484] = 8'd0;
                        text[485] = 8'd0;
                        text[486] = 8'd0;
                        text[487] = 8'd0;
                        text[488] = 8'd0;
                        text[489] = 8'd0;
                        text[490] = 8'd0;
                        text[491] = 8'd0;
                        text[492] = 8'd0;
                        text[493] = 8'd0;
                        text[494] = 8'd0;
                        text[495] = 8'd0;
                        text[496] = 8'd0;
                        text[497] = 8'd0;
                    end else if(text[401] == 8'd71) begin
                        text[401] <= 0;
                        state_R <= 1;
                        ptr <= 32'd401;
                        $display("401 : %d", text[401]);
                        $display("state: %d", state_R);
                        text[480] = 8'd0;
                        text[481] = 8'd0;
                        text[482] = 8'd0;
                        text[483] = 8'd0;
                        text[484] = 8'd0;
                        text[485] = 8'd0;
                        text[486] = 8'd0;
                        text[487] = 8'd0;
                        text[488] = 8'd0;
                        text[489] = 8'd0;
                        text[490] = 8'd0;
                        text[491] = 8'd0;
                        text[492] = 8'd0;
                        text[493] = 8'd0;
                        text[494] = 8'd0;
                        text[495] = 8'd0;
                        text[496] = 8'd0;
                        text[497] = 8'd0;
                    end else if(text[401] == 8'd67) begin
                        text[401] <= 0;
                        state_R <= 4;
                        ptr <= 32'd401;
                        $display("401 : %d", text[401]);
                        $display("state: %d", state_R);
                        text[480] = 8'd0;
                        text[481] = 8'd0;
                        text[482] = 8'd0;
                        text[483] = 8'd0;
                        text[484] = 8'd0;
                        text[485] = 8'd0;
                        text[486] = 8'd0;
                        text[487] = 8'd0;
                        text[488] = 8'd0;
                        text[489] = 8'd0;
                        text[490] = 8'd0;
                        text[491] = 8'd0;
                        text[492] = 8'd0;
                        text[493] = 8'd0;
                        text[494] = 8'd0;
                        text[495] = 8'd0;
                        text[496] = 8'd0;
                        text[497] = 8'd0;
                    end else if(text[401] == 8'd73) begin
                        text[401] <= 0;
                        state_R <= 2;
                        ptr <= 32'd401;
                        $display("401 : %d", text[401]);
                        $display("state: %d", state_R);
                        text[480] = 8'd0;
                        text[481] = 8'd0;
                        text[482] = 8'd0;
                        text[483] = 8'd0;
                        text[484] = 8'd0;
                        text[485] = 8'd0;
                        text[486] = 8'd0;
                        text[487] = 8'd0;
                        text[488] = 8'd0;
                        text[489] = 8'd0;
                        text[490] = 8'd0;
                        text[491] = 8'd0;
                        text[492] = 8'd0;
                        text[493] = 8'd0;
                        text[494] = 8'd0;
                        text[495] = 8'd0;
                        text[496] = 8'd0;
                        text[497] = 8'd0;
                    end else begin// display "Syntax error !!!!!" and clear word typed
                        ptr <= 401;
                        text[480] = 8'd83;
                        text[481] = 8'd121;
                        text[482] = 8'd110;
                        text[483] = 8'd116;
                        text[484] = 8'd97;
                        text[485] = 8'd120;
                        text[486] = 8'd32;
                        text[487] = 8'd101;
                        text[488] = 8'd114;
                        text[489] = 8'd114;
                        text[490] = 8'd111;
                        text[491] = 8'd114;
                        text[492] = 8'd32;
                        text[493] = 8'd33;
                        text[494] = 8'd33;
                        text[495] = 8'd33;
                        text[496] = 8'd33;
                        text[497] = 8'd33;
                        text[401] = 8'd0;
                        text[402] = 8'd0;
                        text[403] = 8'd0;
                        text[404] = 8'd0;
                        text[405] = 8'd0;
                        text[406] = 8'd0;
                        text[407] = 8'd0;
                        text[408] = 8'd0;
                        text[409] = 8'd0;
                        text[410] = 8'd0;
                        text[411] = 8'd0;
                        text[412] = 8'd0;
                        text[413] = 8'd0;
                        text[414] = 8'd0;
                        text[415] = 8'd0;
                        text[416] = 8'd0;
                        text[417] = 8'd0;
                        text[418] = 8'd0;
                        text[419] = 8'd0;
                        text[420] = 8'd0;
                        text[421] = 8'd0;
                        text[422] = 8'd0;
                        text[423] = 8'd0;
                        text[424] = 8'd0;
                        text[425] = 8'd0;
                        text[426] = 8'd0;
                        text[427] = 8'd0;
                        text[428] = 8'd0;
                        text[429] = 8'd0;
                        text[430] = 8'd0;
                        text[431] = 8'd0;
                        text[432] = 8'd0;
                        text[433] = 8'd0;
                        text[434] = 8'd0;
                        text[435] = 8'd0;
                        text[436] = 8'd0;
                        text[437] = 8'd0;
                        text[438] = 8'd0;
                        text[439] = 8'd0;
                        text[440] = 8'd0;
                        text[441] = 8'd0;
                        text[442] = 8'd0;
                        text[443] = 8'd0;
                        text[444] = 8'd0;
                        text[445] = 8'd0;
                        text[446] = 8'd0;
                        text[447] = 8'd0;
                        text[448] = 8'd0;
                        text[449] = 8'd0;
                        text[450] = 8'd0;
                        text[451] = 8'd0;
                        text[452] = 8'd0;
                        text[453] = 8'd0;
                        text[454] = 8'd0;
                        text[455] = 8'd0;
                        text[456] = 8'd0;
                        text[457] = 8'd0;
                        text[458] = 8'd0;
                        text[459] = 8'd0;
                        text[460] = 8'd0;
                        text[461] = 8'd0;
                        text[462] = 8'd0;
                        text[463] = 8'd0;
                        text[464] = 8'd0;
                        text[465] = 8'd0;
                        text[466] = 8'd0;
                        text[467] = 8'd0;
                        text[468] = 8'd0;
                        text[469] = 8'd0;
                        text[470] = 8'd0;
                        text[471] = 8'd0;
                        text[472] = 8'd0;
                        text[473] = 8'd0;
                        text[474] = 8'd0;
                        text[475] = 8'd0;
                        text[476] = 8'd0;
                        text[477] = 8'd0;
                        text[478] = 8'd0;
                        text[479] = 8'd0;
                    end
                end else begin
                    text[ptr] <= ascii_in;
                    if(kbsig[8] == 0 & kbsig[7] == 0 & kbsig[6] == 0 & kbsig[5] == 0 & kbsig[9] == 0)begin
                        ptr <= (ptr < 479) ? ptr + 1 : ptr;
                    end
                end
            end
            else if(kbsig[6] == 1)begin
                ptr <= ((ptr % 80) < 79) ? (ptr + 1) : ptr;
            end
            else if(kbsig[5] == 1)begin
                ptr <= ((ptr % 80) > 0) ? (ptr - 1) : ptr;
            end
            else if(kbsig[9] == 1) begin
                ptr <= (ptr > 401) ? ptr - 1 : ptr;
                if(ptr > 401)begin
                    text[(ptr > 0) ? ptr - 1 : ptr] <= 0;
                end
            end
        end
    end

    get_charpix pix(
        .c(text[80 * (addra / (640 * 16)) + (((addra % (640 * 16)) / 8) % 80)]),
        .x(xw[5:0]),
        .y(yw[5:0]),
        .in_ptr((80 * (addra / (640 * 16)) + (((addra % (640 * 16)) / 8) % 80)) == ptr),
        .is_light(out)
    );

    assign douta = (out == 1) ? 12'b111111111111 : 12'd0; 
endmodule