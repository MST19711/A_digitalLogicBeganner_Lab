`timescale 1ns / 1ps

module mem8b(
   output reg [7:0] dataout,   //???????
   input cs,                   //????????????��????��????��??????????
   input clk,                   //??????
   input we,                   //?��??��????????????????��??????
   input [7:0] datain,        //??????????
   input [15:0] addr         //16��?��????????��????64KB
);

   (* ram_style="block" *) reg [7:0] ram [2**16-1:0];   //????????RAM????��??
    integer i;
    initial
    begin
        for(i = 0; i < 2**16; i = i+1)
        begin
            ram[i] = 8'h00;
        end    
     end 
           
// Add your code here
   
   always @(posedge clk) begin
      dataout <= ram[addr];
   end
   always @(negedge clk) begin
      if (we & cs) ram[addr] <= datain;
   end

endmodule
