`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/09/16 20:18:12
// Design Name: 
// Module Name: regfile32_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module DigitalTimer_tb();
/*
    wire clk;//���ӵ�ʱ�Ӷ˿� CLK100MHZ������ E3
    wire RST;//��λ��ť��������Ч
    wire StartOrPause;//��ʱ����ʼ����ͣ������ 1 �ο�ʼ���ٰ� 1 ����ͣ
    wire ReadPara;//��ȡ���������������ý����󣬵��� 1 �Σ���ȡ����
    wire TimeFormat;//=0 ��ʾ 24 Сʱ�ƣ�=1 ��ʾ 12 Сʱ��
    wire [1:0] mode;//����ѡ��00 ����ʱ�ӣ�01 ����ʱ��10 ��ʱ����11 ��������
    wire [1:0] ParaSelect;// �������ã�00 �ޣ�01 ����������10 ���÷��ӣ�11 ����Сʱ
    wire [1:0] AlarmNo;// ������ţ�0~3
    wire [3:0] data_h;//���ò�����λ��ʹ�� BCD ���ʾ
    wire [3:0] data_l;//���ò�����λ��ʹ�� BCD ���ʾ
    wire Afternoon;//12 Сʱ��ʱ������ʱ�����Ϊ 1
    wire [2:0] TimeKeeper;//������� 3 ɫָʾ��
    wire [2:0] AlarmDisplay;//������� 3 ɫָʾ��
    wire [7:0] segs;//�߶����������ֵ����ʾ����
    wire [7:0] an;//�߶�����ܿ���λ������ʱ���֡���
    DigitalTimer timer_test(
        .clk(clk),//���ӵ�ʱ�Ӷ˿� CLK100MHZ������ E3
        .wire RST(RST),//��λ��ť��������Ч
        .StartOrPause(StartOrPause),//��ʱ����ʼ����ͣ������ 1 �ο�ʼ���ٰ� 1 ����ͣ
        .ReadPara(ReadPara),//��ȡ���������������ý����󣬵��� 1 �Σ���ȡ����
        .TimeFormat(TimeFormat),//=0 ��ʾ 24 Сʱ�ƣ�=1 ��ʾ 12 Сʱ��
        .[1:0] mode(mode),//����ѡ��00 ����ʱ�ӣ�01 ����ʱ��10 ��ʱ����11 ��������
        .[1:0] ParaSelect(ParaSelect),// �������ã�00 �ޣ�01 ����������10 ���÷��ӣ�11 ����Сʱ
        .[1:0] AlarmNo(AlarmNo),// ������ţ�0~3
        .[3:0] data_h(data_h),//���ò�����λ��ʹ�� BCD ���ʾ
        .[3:0] data_l(data_l),//���ò�����λ��ʹ�� BCD ���ʾ
        .Afternoon(Afternoon),//12 Сʱ��ʱ������ʱ�����Ϊ 1
        .[2:0] TimeKeeper(TimeKeeper),//������� 3 ɫָʾ��
        .[2:0] AlarmDisplay(AlarmDisplay),//������� 3 ɫָʾ��
        .[7:0] segs(segs),//�߶����������ֵ����ʾ����
        .[7:0] an(an)//�߶�����ܿ���λ������ʱ���֡���
    );
*/
   

endmodule
